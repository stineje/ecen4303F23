magic
tech scmos
timestamp 1053722803
<< nwell >>
rect -5 48 60 105
<< ntransistor >>
rect 7 6 9 26
rect 23 6 25 26
rect 31 6 33 26
rect 39 6 41 26
rect 47 6 49 26
<< ptransistor >>
rect 7 54 9 94
rect 23 54 25 94
rect 31 54 33 94
rect 39 54 41 94
rect 47 54 49 94
<< ndiffusion >>
rect 6 6 7 26
rect 9 6 10 26
rect 22 6 23 26
rect 25 12 26 26
rect 30 12 31 26
rect 25 6 31 12
rect 33 6 34 26
rect 38 6 39 26
rect 41 23 47 26
rect 41 6 42 23
rect 46 6 47 23
rect 49 23 54 26
rect 49 6 50 23
<< pdiffusion >>
rect 6 54 7 94
rect 9 54 10 94
rect 22 54 23 94
rect 25 88 31 94
rect 25 54 26 88
rect 30 54 31 88
rect 33 54 34 94
rect 38 54 39 94
rect 41 61 42 94
rect 46 61 47 94
rect 41 54 47 61
rect 49 54 50 94
<< ndcontact >>
rect 2 6 6 26
rect 10 6 14 26
rect 18 6 22 26
rect 26 12 30 26
rect 34 6 38 26
rect 42 6 46 23
rect 50 6 54 23
<< pdcontact >>
rect 2 54 6 94
rect 10 54 14 94
rect 18 54 22 94
rect 26 54 30 88
rect 34 54 38 94
rect 42 61 46 94
rect 50 54 54 94
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
rect 46 -2 50 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
rect 46 98 50 102
<< polysilicon >>
rect 7 94 9 96
rect 23 94 25 96
rect 31 94 33 96
rect 39 94 41 96
rect 47 94 49 96
rect 7 51 9 54
rect 23 53 25 54
rect 31 53 33 54
rect 6 49 9 51
rect 12 51 33 53
rect 39 53 41 54
rect 47 53 49 54
rect 39 51 49 53
rect 12 45 14 51
rect 47 37 49 51
rect 7 29 9 33
rect 47 29 49 33
rect 7 27 33 29
rect 7 26 9 27
rect 23 26 25 27
rect 31 26 33 27
rect 39 27 49 29
rect 39 26 41 27
rect 47 26 49 27
rect 7 4 9 6
rect 23 4 25 6
rect 31 4 33 6
rect 39 4 41 6
rect 47 4 49 6
<< polycontact >>
rect 2 47 6 51
rect 10 41 14 45
rect 45 33 49 37
rect 3 29 7 33
<< metal1 >>
rect -2 102 58 103
rect 2 98 14 102
rect 18 98 30 102
rect 34 98 46 102
rect 50 98 58 102
rect -2 97 58 98
rect 2 94 6 97
rect 42 94 46 97
rect 22 91 34 94
rect 38 54 50 58
rect 2 43 6 47
rect 10 45 13 54
rect 26 47 29 54
rect 2 33 5 43
rect 26 43 30 47
rect 2 29 3 33
rect 10 26 13 41
rect 26 26 29 43
rect 49 33 54 37
rect 34 26 54 29
rect 22 6 34 9
rect 51 23 54 26
rect 2 3 6 6
rect 42 3 46 6
rect -2 2 58 3
rect 2 -2 14 2
rect 18 -2 30 2
rect 34 -2 46 2
rect 50 -2 58 2
rect -2 -3 58 -2
<< m1p >>
rect 2 43 6 47
rect 26 43 30 47
rect 50 33 54 37
<< labels >>
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 4 0 4 0 8 gnd
rlabel metal1 52 35 52 35 1 A
rlabel m1p 4 45 4 45 1 EN
rlabel m1p 28 45 28 45 1 Y
<< end >>

VERSION 5.3 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.1 ;

LAYER nwell
  TYPE	MASTERSLICE ;
END nwell

LAYER nactive
  TYPE	MASTERSLICE ;
END nactive

LAYER pactive
  TYPE	MASTERSLICE ;
END pactive

LAYER poly
  TYPE	MASTERSLICE ;
END poly

LAYER cc
  TYPE	CUT ;
  SPACING	0.9 ;
END cc

LAYER metal1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		2.0  ;
  WIDTH		0.6 ;
  SPACING	0.6 ;
  RESISTANCE	RPERSQ 0.07 ;
  CAPACITANCE	CPERSQDIST 3e-5 ;
  CURRENTDEN 0 ;
END metal1

LAYER via
  TYPE	CUT ;
  SPACING	0.6 ;
END via

LAYER metal2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		1.6  ;
  WIDTH		0.6 ;
  SPACING	0.6 ;
  RESISTANCE	RPERSQ 0.07 ;
  CAPACITANCE	CPERSQDIST 1.7e-5 ;
  CURRENTDEN 0 ;
END metal2

LAYER via2
  TYPE	CUT ;
  SPACING	0.6 ;
END via2

LAYER metal3
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		2  ;
  WIDTH		0.6 ;
  SPACING	0.6 ;
  RESISTANCE	RPERSQ 0.07 ;
  CAPACITANCE	CPERSQDIST 7e-6 ;
  CURRENTDEN 0 ;
END metal3

LAYER via3
  TYPE	CUT ;
  SPACING 0.8 ;
END via3

LAYER metal4
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		3.2  ;
  WIDTH		1.2 ;
  SPACING	1.2 ;
  RESISTANCE	RPERSQ 0.04 ;
  CAPACITANCE	CPERSQDIST 4e-6 ;
  CURRENTDEN 0 ;
END metal4

VIA M4_M3 DEFAULT
  LAYER metal3 ;
    RECT -0.400 -0.400 0.400 0.400 ;
  LAYER via3 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER metal4 ;
    RECT -0.600 -0.600 0.600 0.600 ;
END M4_M3

VIA M3_M2 DEFAULT
  LAYER metal2 ;
    RECT -0.400 -0.400 0.400 0.400 ;
  LAYER via2 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER metal3 ;
    RECT -0.400 -0.400 0.400 0.400 ;
END M3_M2

VIA M2_M1 DEFAULT
  LAYER metal1 ;
    RECT -0.400 -0.400 0.400 0.400 ;
  LAYER via ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER metal2 ;
    RECT -0.400 -0.400 0.400 0.400 ;
END M2_M1


VIARULE viagen21 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.6 TO 60 ;
    OVERHANG 0.20 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 0.6 TO 60 ;
    OVERHANG 0.20 ;
    METALOVERHANG 0 ;
  LAYER via ;
    RECT -0.20 -0.20 0.20 0.20 ;
    SPACING 1 BY 1 ;
END viagen21

VIARULE viagen32 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.6 TO 60 ;
    OVERHANG 0.20 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 0.6 TO 60 ;
    OVERHANG 0.20 ;
    METALOVERHANG 0 ;
  LAYER via2 ;
    RECT -0.20 -0.20 0.20 0.20 ;
    SPACING 1 BY 1 ;
END viagen32

VIARULE viagen43 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.6 TO 60 ;
    OVERHANG 0.40 ;
    METALOVERHANG 0 ;
  LAYER metal4 ;
    DIRECTION VERTICAL ;
    WIDTH 0.6 TO 60 ;
    OVERHANG 0.40 ;
    METALOVERHANG 0 ;
  LAYER via3 ;
    RECT -0.20 -0.20 0.20 0.20 ;
    SPACING 1.2 BY 1.2 ;
END viagen43

VIARULE TURN1 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
  LAYER metal1 ;
    DIRECTION VERTICAL ;
END TURN1

VIARULE TURN2 GENERATE
  LAYER metal2 ;
    DIRECTION HORIZONTAL ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
END TURN2

VIARULE TURN3 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
  LAYER metal3 ;
    DIRECTION VERTICAL ;
END TURN3

VIARULE TURN4 GENERATE
  LAYER metal4 ;
    DIRECTION HORIZONTAL ;
  LAYER metal4 ;
    DIRECTION VERTICAL ;
END TURN4

SITE  core
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	1.600 BY 20.000 ;
END  core

SITE  IO
    CLASS	PAD ;
    SYMMETRY	Y ;
    SIZE	90.000 BY 300.000 ;
END  IO

SITE corner
    CLASS 	PAD ;
    SYMMETRY    Y R90 ;
    SIZE 	300.000 BY 300.000 ;
END corner

END LIBRARY

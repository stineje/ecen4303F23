magic
tech sky130A
magscale 1 2
timestamp 1605717589
<< poly >>
rect -16 34 50 44
rect -16 0 0 34
rect 34 0 50 34
rect -16 -10 50 0
<< polycont >>
rect 0 0 34 34
<< locali >>
rect 0 34 34 51
rect 0 -16 34 0
<< end >>

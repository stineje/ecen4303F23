VERSION 5.3 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.075 ;

LAYER nwell
  TYPE	MASTERSLICE ;
END nwell

LAYER nactive
  TYPE	MASTERSLICE ;
END nactive

LAYER pactive
  TYPE	MASTERSLICE ;
END pactive

LAYER poly
  TYPE	MASTERSLICE ;
END poly

LAYER cc
  TYPE	CUT ;
  SPACING	0.450 ;
END cc

LAYER metal1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		1.50  ;
  WIDTH		0.450 ;
  SPACING	0.450 ;
  RESISTANCE	RPERSQ 0.07;
  CAPACITANCE	CPERSQDIST 3.6e-5 ;
  CURRENTDEN 0 ;
END metal1

LAYER via
  TYPE	CUT ;
  SPACING	0.450 ;
END via

LAYER metal2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		1.20  ;
  WIDTH		0.450 ;
  SPACING	0.450 ;
  RESISTANCE	RPERSQ 0.07 ;
  CAPACITANCE	CPERSQDIST 1.6e-5 ;
  CURRENTDEN 0 ;
END metal2

LAYER via2
  TYPE	CUT ;
  SPACING	0.450 ;
END via2

LAYER metal3
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		1.50  ;
  WIDTH		0.450 ;
  SPACING	0.450 ;
  RESISTANCE	RPERSQ 0.07 ;
  CAPACITANCE	CPERSQDIST 1e-5 ;
  CURRENTDEN 0 ;
END metal3

LAYER via3
  TYPE	CUT ;
  SPACING	0.6 ;
END via3

LAYER metal4
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		1.20  ;
  WIDTH		0.450 ;
  SPACING	0.450 ;
  RESISTANCE	RPERSQ 0.07 ;
  CAPACITANCE	CPERSQDIST 5e-6 ;
  CURRENTDEN 0 ;
END metal4

LAYER via4
  TYPE	CUT ;
  SPACING	0.450 ;
END via4

LAYER metal5
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		1.50  ;
  WIDTH		0.60 ;
  SPACING	0.450 ;
  RESISTANCE	RPERSQ 0.02 ;
  CAPACITANCE	CPERSQDIST 4e-6 ;
  CURRENTDEN 0 ;
END metal5

SPACING
END SPACING

VIA M5_M4 DEFAULT
  LAYER metal4 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER via4 ;
    RECT -0.150 -0.150 0.150 0.150 ;
  LAYER metal5 ;
    RECT -0.300 -0.300 0.300 0.300 ;
END M5_M4

VIA M4_M3 DEFAULT
  LAYER metal3 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER via3 ;
    RECT -0.150 -0.150 0.150 0.150 ;
  LAYER metal4 ;
    RECT -0.300 -0.300 0.300 0.300 ;
END M4_M3

VIA M3_M2 DEFAULT
  LAYER metal2 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER via2 ;
    RECT -0.150 -0.150 0.150 0.150 ;
  LAYER metal3 ;
    RECT -0.300 -0.300 0.300 0.300 ;
END M3_M2

VIA M2_M1 DEFAULT
  LAYER metal1 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER via ;
    RECT -0.150 -0.150 0.150 0.150 ;
  LAYER metal2 ;
    RECT -0.300 -0.300 0.300 0.300 ;
END M2_M1

VIARULE viagen21 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.60 TO 60 ;
    OVERHANG 0.150 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 0.6 TO 60 ;
    OVERHANG 0.15 ;
    METALOVERHANG 0 ;
  LAYER via ;
    RECT -0.150 -0.150 0.150 0.150 ;
    SPACING 0.750 BY 0.750 ;
END viagen21

VIARULE viagen32 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.60 TO 60 ;
    OVERHANG 0.15 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 0.6 TO 60 ;
    OVERHANG 0.15 ;
    METALOVERHANG 0 ;
  LAYER via2 ;
    RECT -0.150 -0.150 0.150 0.150 ;
    SPACING 0.750 BY 0.750 ;
END viagen32

VIARULE viagen43 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.60 TO 60 ;
    OVERHANG 0.15 ;
    METALOVERHANG 0 ;
  LAYER metal4 ;
    DIRECTION VERTICAL ;
    WIDTH 0.60 TO 60 ;
    OVERHANG 0.15 ;
    METALOVERHANG 0 ;
  LAYER via3 ;
    RECT -0.150 -0.150 0.150 0.150 ;
    SPACING 0.9 BY 0.9 ;
END viagen43

VIARULE viagen54 GENERATE
  LAYER metal5 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.60 TO 60 ;
    OVERHANG 0.15 ;
    METALOVERHANG 0 ;
  LAYER metal4 ;
    DIRECTION VERTICAL ;
    WIDTH 0.60 TO 60 ;
    OVERHANG 0.150 ;
    METALOVERHANG 0 ;
  LAYER via4 ;
    RECT -0.150 -0.150 0.150 0.150 ;
    SPACING 0.750 BY 0.750 ;
END viagen54


VIARULE TURN1 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
  LAYER metal1 ;
    DIRECTION VERTICAL ;
END TURN1

VIARULE TURN2 GENERATE
  LAYER metal2 ;
    DIRECTION HORIZONTAL ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
END TURN2

VIARULE TURN3 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
  LAYER metal3 ;
    DIRECTION VERTICAL ;
END TURN3

VIARULE TURN4 GENERATE
  LAYER metal4 ;
    DIRECTION HORIZONTAL ;
  LAYER metal4 ;
    DIRECTION VERTICAL ;
END TURN4

VIARULE TURN5 GENERATE
  LAYER metal5 ;
    DIRECTION HORIZONTAL ;
  LAYER metal5 ;
    DIRECTION VERTICAL ;
END TURN5

SITE  core
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	1.200 BY 15.000 ;
END  core

END LIBRARY

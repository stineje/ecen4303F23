magic
tech scmos
timestamp 1053722803
<< nwell >>
rect -5 48 42 105
<< ntransistor >>
rect 7 6 9 16
rect 24 6 26 26
rect 29 6 31 26
<< ptransistor >>
rect 7 74 9 94
rect 24 54 26 94
rect 29 54 31 94
<< ndiffusion >>
rect 6 6 7 16
rect 9 6 10 16
rect 23 6 24 26
rect 26 6 29 26
rect 31 6 32 26
<< pdiffusion >>
rect 6 74 7 94
rect 9 74 10 94
rect 23 54 24 94
rect 26 54 29 94
rect 31 54 32 94
<< ndcontact >>
rect 2 6 6 16
rect 10 6 14 16
rect 19 6 23 26
rect 32 6 36 26
<< pdcontact >>
rect 2 74 6 94
rect 10 74 14 94
rect 19 54 23 94
rect 32 54 36 94
<< psubstratepcontact >>
rect -2 -2 2 2
rect 22 -2 26 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 22 98 26 102
<< polysilicon >>
rect 7 94 9 96
rect 24 94 26 96
rect 29 94 31 96
rect 7 67 9 74
rect 7 29 9 63
rect 24 35 26 54
rect 17 33 26 35
rect 29 37 31 54
rect 29 33 30 37
rect 7 27 26 29
rect 7 16 9 27
rect 24 26 26 27
rect 29 26 31 33
rect 7 4 9 6
rect 24 4 26 6
rect 29 4 31 6
<< polycontact >>
rect 6 63 10 67
rect 13 33 17 37
rect 30 33 34 37
<< metal1 >>
rect -2 102 42 103
rect 2 98 22 102
rect 26 98 42 102
rect -2 97 42 98
rect 2 94 6 97
rect 32 94 36 97
rect 14 74 16 77
rect 2 63 6 67
rect 13 53 16 74
rect 12 50 16 53
rect 12 40 15 50
rect 20 47 23 54
rect 18 43 23 47
rect 12 37 16 40
rect 13 16 16 33
rect 20 26 23 43
rect 34 33 38 37
rect 14 12 16 16
rect 2 3 6 6
rect 32 3 36 6
rect -2 2 42 3
rect 2 -2 22 2
rect 26 -2 42 2
rect -2 -3 42 -2
<< m1p >>
rect 2 63 6 67
rect 18 43 22 47
rect 34 33 38 37
<< labels >>
<< end >>

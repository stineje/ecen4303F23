magic
tech scmos
timestamp 1053722803
<< nwell >>
rect -9 48 28 105
<< ntransistor >>
rect 7 6 9 26
rect 15 6 17 26
<< ptransistor >>
rect 7 54 9 94
rect 15 54 17 94
<< ndiffusion >>
rect 6 6 7 26
rect 9 6 10 26
rect 14 6 15 26
rect 17 6 18 26
<< pdiffusion >>
rect 6 54 7 94
rect 9 54 10 94
rect 14 54 15 94
rect 17 54 18 94
<< ndcontact >>
rect 2 6 6 26
rect 10 6 14 26
rect 18 6 22 26
<< pdcontact >>
rect 2 54 6 94
rect 10 54 14 94
rect 18 54 22 94
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 7 53 9 54
rect 15 53 17 54
rect 7 51 17 53
rect 7 33 9 51
rect 6 30 9 33
rect 6 29 17 30
rect 7 28 17 29
rect 7 26 9 28
rect 15 26 17 28
rect 7 4 9 6
rect 15 4 17 6
<< polycontact >>
rect 2 29 6 33
<< metal1 >>
rect -2 102 26 103
rect 2 98 14 102
rect 18 98 26 102
rect -2 97 26 98
rect 2 94 6 97
rect 18 94 22 97
rect 2 33 6 37
rect 10 26 14 54
rect 2 3 6 6
rect 18 3 22 6
rect -2 2 26 3
rect 2 -2 14 2
rect 18 -2 26 2
rect -2 -3 26 -2
<< m1p >>
rect 10 43 14 47
rect 2 33 6 37
<< labels >>
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 4 0 4 0 8 gnd
rlabel m1p 12 45 12 45 6 Y
rlabel m1p 4 35 4 35 6 A
<< end >>

magic
tech scmos
timestamp 1053722803
<< nwell >>
rect -9 48 37 105
<< ntransistor >>
rect 7 6 9 21
rect 15 6 17 26
rect 23 6 25 26
<< ptransistor >>
rect 7 64 9 94
rect 15 54 17 94
rect 23 54 25 94
<< ndiffusion >>
rect 6 6 7 21
rect 9 6 10 21
rect 14 6 15 26
rect 17 6 18 26
rect 22 6 23 26
rect 25 6 26 26
<< pdiffusion >>
rect 6 64 7 94
rect 9 64 10 94
rect 14 60 15 94
rect 10 54 15 60
rect 17 54 18 94
rect 22 54 23 94
rect 25 54 26 94
<< ndcontact >>
rect 2 6 6 21
rect 10 6 14 26
rect 18 6 22 26
rect 26 6 30 26
<< pdcontact >>
rect 2 64 6 94
rect 10 60 14 94
rect 18 54 22 94
rect 26 54 30 94
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 7 21 9 64
rect 15 53 17 54
rect 23 53 25 54
rect 15 51 25 53
rect 15 44 17 51
rect 15 29 17 40
rect 15 27 25 29
rect 15 26 17 27
rect 23 26 25 27
rect 7 4 9 6
rect 15 4 17 6
rect 23 4 25 6
<< polycontact >>
rect 3 39 7 43
rect 13 40 17 44
<< metal1 >>
rect -2 102 34 103
rect 2 98 14 102
rect 18 98 34 102
rect -2 97 34 98
rect 10 94 14 97
rect 26 94 30 97
rect 2 57 6 64
rect 2 54 15 57
rect 22 54 23 59
rect 2 43 7 47
rect 12 44 15 54
rect 12 40 13 44
rect 12 32 15 40
rect 20 37 23 54
rect 18 33 23 37
rect 2 29 15 32
rect 2 21 6 29
rect 20 26 23 33
rect 22 23 23 26
rect 10 3 14 6
rect 26 3 30 6
rect -2 2 34 3
rect 2 -2 14 2
rect 18 -2 34 2
rect -2 -3 34 -2
<< m1p >>
rect 2 43 6 47
rect 18 33 22 37
<< labels >>
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1600264764
<< nwell >>
rect -100 161 136 448
<< nmos >>
rect 0 -41 30 43
<< pmos >>
rect 0 197 30 281
<< ndiff >>
rect -73 3 0 43
rect -73 -33 -48 3
rect -14 -33 0 3
rect -73 -41 0 -33
rect 30 3 91 43
rect 30 -33 41 3
rect 75 -33 91 3
rect 30 -41 91 -33
<< pdiff >>
rect -57 273 0 281
rect -57 237 -45 273
rect -11 237 0 273
rect -57 197 0 237
rect 30 273 87 281
rect 30 237 41 273
rect 75 237 87 273
rect 30 197 87 237
<< ndiffc >>
rect -48 -33 -14 3
rect 41 -33 75 3
<< pdiffc >>
rect -45 237 -11 273
rect 41 237 75 273
<< psubdiff >>
rect -17 -142 7 -106
rect 43 -142 67 -106
<< nsubdiff >>
rect -22 346 2 382
rect 38 346 62 382
<< psubdiffcont >>
rect 7 -142 43 -106
<< nsubdiffcont >>
rect 2 346 38 382
<< poly >>
rect 0 281 30 323
rect 0 150 30 197
rect -64 134 30 150
rect -64 91 -48 134
rect 0 91 30 134
rect -64 75 30 91
rect 0 43 30 75
rect 0 -73 30 -41
<< polycont >>
rect -48 91 0 134
<< locali >>
rect -113 382 166 394
rect -113 346 2 382
rect 38 346 166 382
rect -113 325 166 346
rect -45 273 -11 325
rect -45 221 -11 237
rect 41 273 75 290
rect -48 134 0 150
rect -48 75 0 91
rect -48 3 -14 19
rect -48 -90 -14 -33
rect 41 3 75 237
rect 41 -53 75 -33
rect -122 -106 157 -90
rect -122 -142 7 -106
rect 43 -142 157 -106
rect -122 -159 157 -142
<< labels >>
rlabel locali 62 135 62 135 1 Y
port 1 n
rlabel locali -24 113 -24 113 1 A
port 2 n
rlabel locali 25 -124 25 -124 1 GND
rlabel locali 17 364 17 364 1 VDD
<< end >>

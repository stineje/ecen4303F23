magic
tech scmos
timestamp 1053022145
<< nwell >>
rect -7 48 68 105
<< ntransistor >>
rect 15 6 17 16
rect 23 6 25 16
rect 31 6 33 16
<< ptransistor >>
rect 7 64 9 94
rect 15 64 17 94
rect 23 64 25 94
rect 31 64 33 94
rect 47 60 49 90
rect 55 60 57 90
<< ndiffusion >>
rect 14 6 15 16
rect 17 6 18 16
rect 22 6 23 16
rect 25 14 31 16
rect 25 6 26 14
rect 30 6 31 14
rect 33 6 34 16
<< pdiffusion >>
rect 6 64 7 94
rect 9 64 10 94
rect 14 64 15 94
rect 17 64 18 94
rect 22 64 23 94
rect 25 88 31 94
rect 25 64 26 88
rect 30 64 31 88
rect 33 65 34 94
rect 33 64 36 65
rect 46 60 47 90
rect 49 88 55 90
rect 49 60 50 88
rect 54 60 55 88
rect 57 60 58 90
<< ndcontact >>
rect 10 6 14 16
rect 18 6 22 16
rect 26 6 30 14
rect 34 6 38 16
<< pdcontact >>
rect 2 64 6 94
rect 10 64 14 94
rect 18 64 22 94
rect 26 64 30 88
rect 34 65 38 94
rect 42 60 46 90
rect 50 60 54 88
rect 58 60 62 90
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
rect 46 -2 50 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
rect 46 98 50 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 31 94 33 96
rect 47 90 49 92
rect 55 90 57 92
rect 7 63 9 64
rect 15 63 17 64
rect 23 63 25 64
rect 31 63 33 64
rect 7 61 17 63
rect 15 27 17 61
rect 22 61 33 63
rect 22 37 24 61
rect 47 59 49 60
rect 55 59 57 60
rect 47 57 57 59
rect 47 56 49 57
rect 31 54 49 56
rect 31 47 33 54
rect 15 16 17 23
rect 23 16 25 33
rect 31 16 33 43
rect 15 4 17 6
rect 23 4 25 6
rect 31 4 33 6
<< polycontact >>
rect 30 43 34 47
rect 22 33 26 37
rect 15 23 19 27
<< metal1 >>
rect -2 102 66 103
rect 2 98 14 102
rect 18 98 30 102
rect 34 98 46 102
rect 50 98 66 102
rect -2 97 66 98
rect 10 94 14 97
rect 22 91 34 94
rect 43 91 61 94
rect 43 90 46 91
rect 3 61 6 64
rect 18 61 21 64
rect 3 58 21 61
rect 27 62 30 64
rect 27 60 42 62
rect 58 90 61 91
rect 27 59 45 60
rect 50 57 53 60
rect 50 56 54 57
rect 37 53 54 56
rect 26 43 30 47
rect 18 33 22 37
rect 10 23 15 27
rect 37 20 40 53
rect 20 17 40 20
rect 20 16 23 17
rect 22 13 23 16
rect 34 16 40 17
rect 10 3 14 6
rect 26 3 30 6
rect -2 2 66 3
rect 2 -2 14 2
rect 18 -2 30 2
rect 34 -2 46 2
rect 50 -2 66 2
rect -2 -3 66 -2
<< m1p >>
rect 50 53 54 57
rect 26 43 30 47
rect 18 33 22 37
rect 10 23 14 27
<< labels >>
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 4 0 4 0 8 gnd
rlabel m1p 20 35 20 35 6 B
rlabel m1p 28 45 28 45 6 C
rlabel m1p 12 25 12 25 6 A
rlabel m1p 52 55 52 55 6 Y
<< end >>

magic
tech scmos
timestamp 1091055042
<< nwell >>
rect 30 1110 420 1500
rect 229 416 271 478
rect 34 409 271 416
rect 34 394 44 409
rect 228 394 271 409
rect 365 411 425 416
rect 365 406 409 411
rect 400 394 409 406
<< pwell >>
rect 224 597 435 599
rect 224 579 226 597
rect 15 576 226 579
rect 269 585 327 597
rect 15 574 231 576
rect 229 535 231 574
rect 269 535 271 585
rect 325 576 327 585
rect 423 576 435 577
rect 325 575 435 576
rect 325 574 425 575
<< hvnwell >>
rect 17 637 433 993
rect -3 478 453 493
rect -3 416 229 478
rect 271 416 453 478
rect -3 394 34 416
rect 44 394 228 409
rect 271 406 365 416
rect 425 411 453 416
rect 271 394 400 406
rect 409 394 453 411
rect -3 378 453 394
rect -3 11 11 378
rect 439 11 453 378
rect -3 -3 453 11
<< hvpwell >>
rect -3 996 453 1013
rect -3 634 14 996
rect 436 634 453 996
rect -3 599 453 634
rect -3 579 224 599
rect 435 597 453 599
rect -3 574 15 579
rect -3 535 229 574
rect -3 534 231 535
rect 271 574 325 585
rect 436 577 453 597
rect 435 575 453 577
rect 425 574 453 575
rect 271 535 453 574
rect 269 534 453 535
rect -3 517 453 534
rect 11 11 439 378
<< hvntransistor >>
rect 20 540 23 570
rect 29 540 32 570
rect 46 540 49 570
rect 55 540 58 570
rect 64 540 67 570
rect 73 540 76 570
rect 82 540 85 570
rect 91 540 94 570
rect 100 540 103 570
rect 109 540 112 570
rect 118 540 121 570
rect 127 540 130 570
rect 136 540 139 570
rect 145 540 148 570
rect 154 540 157 570
rect 163 540 166 570
rect 180 540 183 570
rect 189 540 192 570
rect 207 540 210 570
rect 216 540 219 570
rect 326 540 329 570
rect 335 540 338 570
rect 344 540 347 570
rect 353 540 356 570
rect 362 540 365 570
rect 371 540 374 570
rect 380 540 383 570
rect 389 540 392 570
rect 398 540 401 570
rect 407 540 410 570
rect 416 540 419 570
rect 425 540 428 570
rect 38 345 213 348
rect 237 345 412 348
rect 38 284 213 287
rect 237 284 412 287
rect 38 263 213 266
rect 237 263 412 266
rect 38 203 213 206
rect 38 182 213 185
rect 237 203 412 206
rect 237 182 412 185
rect 38 122 213 125
rect 237 122 412 125
rect 38 101 213 104
rect 237 101 412 104
rect 38 41 213 44
rect 237 41 412 44
<< hvptransistor >>
rect 38 965 213 968
rect 237 965 412 968
rect 38 904 213 907
rect 237 904 412 907
rect 38 883 213 886
rect 237 883 412 886
rect 38 823 213 826
rect 237 823 412 826
rect 38 802 213 805
rect 237 802 412 805
rect 38 742 213 745
rect 237 742 412 745
rect 38 721 213 724
rect 237 721 412 724
rect 38 661 213 664
rect 237 661 412 664
rect 20 420 23 472
rect 29 420 32 472
rect 46 420 49 472
rect 55 420 58 472
rect 64 420 67 472
rect 73 420 76 472
rect 82 420 85 472
rect 91 420 94 472
rect 100 420 103 472
rect 109 420 112 472
rect 118 420 121 472
rect 127 420 130 472
rect 136 420 139 472
rect 145 420 148 472
rect 154 420 157 472
rect 163 420 166 472
rect 181 420 184 472
rect 190 420 193 472
rect 208 420 211 472
rect 217 420 220 472
rect 326 420 329 472
rect 335 420 338 472
rect 344 420 347 472
rect 353 420 356 472
rect 362 420 365 472
rect 371 420 374 472
rect 380 420 383 472
rect 389 420 392 472
rect 398 420 401 472
rect 407 420 410 472
rect 416 420 419 472
rect 425 420 428 472
<< hvndiffusion >>
rect 11 584 19 618
rect 23 614 39 618
rect 173 614 437 618
rect 23 613 437 614
rect 23 609 275 613
rect 434 609 437 613
rect 23 608 437 609
rect 23 604 39 608
rect 173 604 437 608
rect 23 603 437 604
rect 23 598 220 603
rect 23 594 39 598
rect 173 594 220 598
rect 23 588 220 594
rect 23 584 39 588
rect 173 584 220 588
rect 11 583 220 584
rect 275 575 321 581
rect 275 571 278 575
rect 317 571 321 575
rect 275 570 321 571
rect 429 570 437 571
rect 19 546 20 570
rect 15 540 20 546
rect 23 569 29 570
rect 23 560 24 569
rect 28 560 29 569
rect 23 555 29 560
rect 23 551 24 555
rect 28 551 29 555
rect 23 545 29 551
rect 23 541 24 545
rect 28 541 29 545
rect 23 540 29 541
rect 32 541 33 570
rect 32 540 37 541
rect 45 541 46 570
rect 41 540 46 541
rect 49 564 55 570
rect 49 560 50 564
rect 54 560 55 564
rect 49 555 55 560
rect 49 551 50 555
rect 54 551 55 555
rect 49 545 55 551
rect 49 541 50 545
rect 54 541 55 545
rect 49 540 55 541
rect 58 541 59 570
rect 63 541 64 570
rect 58 540 64 541
rect 67 564 73 570
rect 67 560 68 564
rect 72 560 73 564
rect 67 555 73 560
rect 67 551 68 555
rect 72 551 73 555
rect 67 545 73 551
rect 67 541 68 545
rect 72 541 73 545
rect 67 540 73 541
rect 76 541 77 570
rect 81 541 82 570
rect 76 540 82 541
rect 85 564 91 570
rect 85 560 86 564
rect 90 560 91 564
rect 85 555 91 560
rect 85 551 86 555
rect 90 551 91 555
rect 85 545 91 551
rect 85 541 86 545
rect 90 541 91 545
rect 85 540 91 541
rect 94 541 95 570
rect 99 541 100 570
rect 94 540 100 541
rect 103 564 109 570
rect 103 560 104 564
rect 108 560 109 564
rect 103 555 109 560
rect 103 551 104 555
rect 108 551 109 555
rect 103 545 109 551
rect 103 541 104 545
rect 108 541 109 545
rect 103 540 109 541
rect 112 541 113 570
rect 117 541 118 570
rect 112 540 118 541
rect 121 564 127 570
rect 121 560 122 564
rect 126 560 127 564
rect 121 555 127 560
rect 121 551 122 555
rect 126 551 127 555
rect 121 545 127 551
rect 121 541 122 545
rect 126 541 127 545
rect 121 540 127 541
rect 130 569 136 570
rect 130 550 131 569
rect 135 550 136 569
rect 130 540 136 550
rect 139 541 140 570
rect 144 541 145 570
rect 139 540 145 541
rect 148 564 154 570
rect 148 550 149 564
rect 153 550 154 564
rect 148 545 154 550
rect 148 541 149 545
rect 153 541 154 545
rect 148 540 154 541
rect 157 546 158 570
rect 162 546 163 570
rect 157 540 163 546
rect 166 541 167 570
rect 166 540 171 541
rect 179 541 180 570
rect 175 540 180 541
rect 183 569 189 570
rect 183 560 184 569
rect 188 560 189 569
rect 183 555 189 560
rect 183 551 184 555
rect 188 551 189 555
rect 183 545 189 551
rect 183 541 184 545
rect 188 541 189 545
rect 183 540 189 541
rect 192 546 194 570
rect 192 540 198 546
rect 206 541 207 570
rect 202 540 207 541
rect 210 569 216 570
rect 210 560 211 569
rect 215 560 216 569
rect 210 555 216 560
rect 210 551 211 555
rect 215 551 216 555
rect 210 545 216 551
rect 210 541 211 545
rect 215 541 216 545
rect 210 540 216 541
rect 219 546 221 570
rect 219 540 225 546
rect 275 565 326 570
rect 275 561 276 565
rect 325 561 326 565
rect 275 555 326 561
rect 275 551 276 555
rect 325 551 326 555
rect 275 545 326 551
rect 275 541 276 545
rect 325 541 326 545
rect 275 540 326 541
rect 329 541 330 570
rect 334 541 335 570
rect 329 540 335 541
rect 338 564 344 570
rect 338 560 339 564
rect 343 560 344 564
rect 338 555 344 560
rect 338 551 339 555
rect 343 551 344 555
rect 338 545 344 551
rect 338 541 339 545
rect 343 541 344 545
rect 338 540 344 541
rect 347 541 348 570
rect 352 541 353 570
rect 347 540 353 541
rect 356 564 362 570
rect 356 560 357 564
rect 361 560 362 564
rect 356 555 362 560
rect 356 551 357 555
rect 361 551 362 555
rect 356 545 362 551
rect 356 541 357 545
rect 361 541 362 545
rect 356 540 362 541
rect 365 541 366 570
rect 370 541 371 570
rect 365 540 371 541
rect 374 569 380 570
rect 374 560 375 569
rect 379 560 380 569
rect 374 555 380 560
rect 374 551 375 555
rect 379 551 380 555
rect 374 545 380 551
rect 374 541 375 545
rect 379 541 380 545
rect 374 540 380 541
rect 383 541 384 570
rect 388 541 389 570
rect 383 540 389 541
rect 392 564 398 570
rect 392 560 393 564
rect 397 560 398 564
rect 392 555 398 560
rect 392 551 393 555
rect 397 551 398 555
rect 392 545 398 551
rect 392 541 393 545
rect 397 541 398 545
rect 392 540 398 541
rect 401 541 402 570
rect 406 541 407 570
rect 401 540 407 541
rect 410 564 416 570
rect 410 560 411 564
rect 415 560 416 564
rect 410 555 416 560
rect 410 551 411 555
rect 415 551 416 555
rect 410 545 416 551
rect 410 541 411 545
rect 415 541 416 545
rect 410 540 416 541
rect 419 541 420 570
rect 424 541 425 570
rect 419 540 425 541
rect 428 569 437 570
rect 428 560 429 569
rect 433 560 437 569
rect 428 555 437 560
rect 428 551 429 555
rect 433 551 437 555
rect 428 545 437 551
rect 428 541 429 545
rect 433 541 437 545
rect 428 540 437 541
rect 50 533 54 540
rect 68 533 72 540
rect 86 533 90 540
rect 122 533 126 540
rect 275 533 325 540
rect 339 533 343 540
rect 357 533 361 540
rect 375 533 379 540
rect 393 533 397 540
rect 411 533 415 540
rect 429 533 437 540
rect 38 356 213 357
rect 38 352 50 356
rect 174 352 213 356
rect 38 348 213 352
rect 38 321 213 345
rect 38 317 56 321
rect 195 317 213 321
rect 38 315 213 317
rect 38 311 56 315
rect 195 311 213 315
rect 38 287 213 311
rect 237 356 412 357
rect 237 352 278 356
rect 397 352 412 356
rect 237 348 412 352
rect 38 280 213 284
rect 38 276 51 280
rect 185 276 213 280
rect 38 274 213 276
rect 38 270 51 274
rect 185 270 213 274
rect 38 266 213 270
rect 237 321 412 345
rect 237 317 255 321
rect 394 317 412 321
rect 237 315 412 317
rect 237 311 255 315
rect 394 311 412 315
rect 237 287 412 311
rect 237 280 412 284
rect 237 276 265 280
rect 399 276 412 280
rect 237 274 412 276
rect 237 270 265 274
rect 399 270 412 274
rect 237 266 412 270
rect 38 239 213 263
rect 38 230 56 239
rect 195 230 213 239
rect 38 206 213 230
rect 38 199 213 203
rect 38 195 51 199
rect 185 195 213 199
rect 38 193 213 195
rect 38 189 51 193
rect 185 189 213 193
rect 38 185 213 189
rect 38 158 213 182
rect 38 149 56 158
rect 195 149 213 158
rect 38 125 213 149
rect 237 239 412 263
rect 237 230 255 239
rect 394 230 412 239
rect 237 206 412 230
rect 237 199 412 203
rect 237 195 265 199
rect 399 195 412 199
rect 237 193 412 195
rect 237 189 265 193
rect 399 189 412 193
rect 237 185 412 189
rect 237 158 412 182
rect 237 149 255 158
rect 394 149 412 158
rect 237 125 412 149
rect 38 118 213 122
rect 38 114 51 118
rect 185 114 213 118
rect 38 112 213 114
rect 38 108 51 112
rect 185 108 213 112
rect 38 104 213 108
rect 38 77 213 101
rect 38 68 56 77
rect 195 68 213 77
rect 38 44 213 68
rect 237 118 412 122
rect 237 114 265 118
rect 399 114 412 118
rect 237 112 412 114
rect 237 108 265 112
rect 399 108 412 112
rect 237 104 412 108
rect 38 37 213 41
rect 38 33 51 37
rect 170 33 213 37
rect 38 32 213 33
rect 237 77 412 101
rect 237 68 255 77
rect 394 68 412 77
rect 237 44 412 68
rect 237 37 412 41
rect 237 33 280 37
rect 399 33 412 37
rect 237 32 412 33
<< hvpdiffusion >>
rect 38 976 213 977
rect 38 972 41 976
rect 170 972 213 976
rect 38 968 213 972
rect 38 941 213 965
rect 38 937 61 941
rect 195 937 213 941
rect 38 935 213 937
rect 38 931 61 935
rect 195 931 213 935
rect 38 907 213 931
rect 237 976 412 977
rect 237 972 280 976
rect 409 972 412 976
rect 237 968 412 972
rect 237 941 412 965
rect 237 937 255 941
rect 389 937 412 941
rect 237 935 412 937
rect 237 931 255 935
rect 389 931 412 935
rect 237 907 412 931
rect 38 900 213 904
rect 38 896 46 900
rect 190 896 213 900
rect 38 894 213 896
rect 38 890 46 894
rect 190 890 213 894
rect 38 886 213 890
rect 237 900 412 904
rect 237 896 260 900
rect 404 896 412 900
rect 237 894 412 896
rect 237 890 260 894
rect 404 890 412 894
rect 237 886 412 890
rect 38 859 213 883
rect 38 850 61 859
rect 195 850 213 859
rect 38 826 213 850
rect 237 859 412 883
rect 237 850 255 859
rect 389 850 412 859
rect 237 826 412 850
rect 38 819 213 823
rect 38 815 46 819
rect 190 815 213 819
rect 38 813 213 815
rect 38 809 46 813
rect 190 809 213 813
rect 38 805 213 809
rect 38 778 213 802
rect 38 769 61 778
rect 195 769 213 778
rect 38 745 213 769
rect 237 819 412 823
rect 237 815 255 819
rect 404 815 412 819
rect 237 813 412 815
rect 237 809 260 813
rect 404 809 412 813
rect 237 805 412 809
rect 38 738 213 742
rect 38 734 46 738
rect 190 734 213 738
rect 38 732 213 734
rect 38 728 46 732
rect 190 728 213 732
rect 38 724 213 728
rect 237 778 412 802
rect 237 769 255 778
rect 389 769 412 778
rect 237 745 412 769
rect 237 738 412 742
rect 237 734 260 738
rect 404 734 412 738
rect 237 732 412 734
rect 237 728 260 732
rect 404 728 412 732
rect 237 724 412 728
rect 38 697 213 721
rect 38 688 61 697
rect 195 688 213 697
rect 38 664 213 688
rect 38 657 213 661
rect 38 653 41 657
rect 170 653 213 657
rect 38 652 213 653
rect 237 697 412 721
rect 237 688 255 697
rect 389 688 412 697
rect 237 664 412 688
rect 237 657 412 661
rect 237 653 280 657
rect 409 653 412 657
rect 237 652 412 653
rect 50 472 54 480
rect 68 472 72 480
rect 86 472 90 480
rect 122 472 126 480
rect 275 477 325 478
rect 275 473 276 477
rect 275 472 325 473
rect 429 472 440 480
rect 15 465 20 472
rect 19 421 20 465
rect 15 420 20 421
rect 23 466 29 472
rect 23 462 24 466
rect 28 462 29 466
rect 23 456 29 462
rect 23 452 24 456
rect 28 452 29 456
rect 23 446 29 452
rect 23 442 24 446
rect 28 442 29 446
rect 23 436 29 442
rect 23 432 24 436
rect 28 432 29 436
rect 23 420 29 432
rect 32 471 37 472
rect 32 422 33 471
rect 32 420 37 422
rect 41 471 46 472
rect 45 422 46 471
rect 41 420 46 422
rect 49 466 55 472
rect 49 462 50 466
rect 54 462 55 466
rect 49 456 55 462
rect 49 452 50 456
rect 54 452 55 456
rect 49 446 55 452
rect 49 442 50 446
rect 54 442 55 446
rect 49 436 55 442
rect 49 432 50 436
rect 54 432 55 436
rect 49 420 55 432
rect 58 471 64 472
rect 58 422 59 471
rect 63 422 64 471
rect 58 420 64 422
rect 67 466 73 472
rect 67 462 68 466
rect 72 462 73 466
rect 67 456 73 462
rect 67 452 68 456
rect 72 452 73 456
rect 67 446 73 452
rect 67 442 68 446
rect 72 442 73 446
rect 67 436 73 442
rect 67 432 68 436
rect 72 432 73 436
rect 67 420 73 432
rect 76 471 82 472
rect 76 422 77 471
rect 81 422 82 471
rect 76 420 82 422
rect 85 466 91 472
rect 85 462 86 466
rect 90 462 91 466
rect 85 456 91 462
rect 85 452 86 456
rect 90 452 91 456
rect 85 446 91 452
rect 85 442 86 446
rect 90 442 91 446
rect 85 436 91 442
rect 85 432 86 436
rect 90 432 91 436
rect 85 420 91 432
rect 94 471 100 472
rect 94 422 95 471
rect 99 422 100 471
rect 94 420 100 422
rect 103 466 109 472
rect 103 462 104 466
rect 108 462 109 466
rect 103 456 109 462
rect 103 452 104 456
rect 108 452 109 456
rect 103 446 109 452
rect 103 442 104 446
rect 108 442 109 446
rect 103 436 109 442
rect 103 432 104 436
rect 108 432 109 436
rect 103 420 109 432
rect 112 471 118 472
rect 112 422 113 471
rect 117 422 118 471
rect 112 420 118 422
rect 121 466 127 472
rect 121 462 122 466
rect 126 462 127 466
rect 121 456 127 462
rect 121 452 122 456
rect 126 452 127 456
rect 121 446 127 452
rect 121 442 122 446
rect 126 442 127 446
rect 121 436 127 442
rect 121 432 122 436
rect 126 432 127 436
rect 121 420 127 432
rect 130 471 136 472
rect 130 422 131 471
rect 135 422 136 471
rect 130 420 136 422
rect 139 466 145 472
rect 139 422 140 466
rect 144 422 145 466
rect 139 420 145 422
rect 148 470 154 472
rect 148 466 149 470
rect 153 466 154 470
rect 148 461 154 466
rect 148 427 149 461
rect 153 427 154 461
rect 148 420 154 427
rect 157 471 163 472
rect 157 422 158 471
rect 162 422 163 471
rect 157 420 163 422
rect 166 461 172 472
rect 166 422 167 461
rect 171 422 172 461
rect 166 420 172 422
rect 175 471 181 472
rect 175 422 176 471
rect 180 422 181 471
rect 175 420 181 422
rect 184 466 190 472
rect 184 462 185 466
rect 189 462 190 466
rect 184 456 190 462
rect 184 452 185 456
rect 189 452 190 456
rect 184 446 190 452
rect 184 442 185 446
rect 189 442 190 446
rect 184 436 190 442
rect 184 432 185 436
rect 189 432 190 436
rect 184 420 190 432
rect 193 466 198 472
rect 193 422 194 466
rect 193 420 198 422
rect 202 471 208 472
rect 202 422 203 471
rect 207 422 208 471
rect 202 420 208 422
rect 211 466 217 472
rect 211 462 212 466
rect 216 462 217 466
rect 211 456 217 462
rect 211 452 212 456
rect 216 452 217 456
rect 211 446 217 452
rect 211 442 212 446
rect 216 442 217 446
rect 211 436 217 442
rect 211 432 212 436
rect 216 432 217 436
rect 211 420 217 432
rect 220 466 225 472
rect 220 422 221 466
rect 220 420 225 422
rect 275 467 326 472
rect 275 463 276 467
rect 325 463 326 467
rect 275 457 326 463
rect 275 453 276 457
rect 325 453 326 457
rect 275 447 326 453
rect 275 443 276 447
rect 325 443 326 447
rect 275 437 326 443
rect 275 433 276 437
rect 325 433 326 437
rect 275 427 326 433
rect 275 423 276 427
rect 325 423 326 427
rect 275 420 326 423
rect 329 471 335 472
rect 329 422 330 471
rect 334 422 335 471
rect 329 420 335 422
rect 338 466 344 472
rect 338 462 339 466
rect 343 462 344 466
rect 338 456 344 462
rect 338 452 339 456
rect 343 452 344 456
rect 338 445 344 452
rect 338 441 339 445
rect 343 441 344 445
rect 338 436 344 441
rect 338 432 339 436
rect 343 432 344 436
rect 338 420 344 432
rect 347 471 353 472
rect 347 427 348 471
rect 352 427 353 471
rect 347 420 353 427
rect 356 466 362 472
rect 356 462 357 466
rect 361 462 362 466
rect 356 456 362 462
rect 356 452 357 456
rect 361 452 362 456
rect 356 445 362 452
rect 356 441 357 445
rect 361 441 362 445
rect 356 436 362 441
rect 356 432 357 436
rect 361 432 362 436
rect 356 420 362 432
rect 365 471 371 472
rect 365 422 366 471
rect 370 422 371 471
rect 365 420 371 422
rect 374 466 380 472
rect 374 462 375 466
rect 379 462 380 466
rect 374 456 380 462
rect 374 452 375 456
rect 379 452 380 456
rect 374 445 380 452
rect 374 441 375 445
rect 379 441 380 445
rect 374 436 380 441
rect 374 432 375 436
rect 379 432 380 436
rect 374 420 380 432
rect 383 471 389 472
rect 383 422 384 471
rect 388 422 389 471
rect 383 420 389 422
rect 392 466 398 472
rect 392 462 393 466
rect 397 462 398 466
rect 392 456 398 462
rect 392 452 393 456
rect 397 452 398 456
rect 392 445 398 452
rect 392 441 393 445
rect 397 441 398 445
rect 392 436 398 441
rect 392 432 393 436
rect 397 432 398 436
rect 392 420 398 432
rect 401 471 407 472
rect 401 422 402 471
rect 406 422 407 471
rect 401 420 407 422
rect 410 470 416 472
rect 410 466 411 470
rect 415 466 416 470
rect 410 461 416 466
rect 410 457 411 461
rect 415 457 416 461
rect 410 451 416 457
rect 410 447 411 451
rect 415 447 416 451
rect 410 441 416 447
rect 410 437 411 441
rect 415 437 416 441
rect 410 431 416 437
rect 410 427 411 431
rect 415 427 416 431
rect 410 420 416 427
rect 419 471 425 472
rect 419 422 420 471
rect 424 422 425 471
rect 419 420 425 422
rect 428 420 429 472
rect 275 417 325 420
rect 19 406 30 411
rect 275 413 276 417
rect 325 413 326 416
rect 19 402 20 406
rect 29 402 30 406
rect 275 408 326 413
rect 433 408 440 472
rect 275 407 361 408
rect 429 407 440 408
rect 19 396 30 402
rect 19 392 20 396
rect 29 392 30 396
rect 48 397 224 405
rect 48 393 49 397
rect 223 393 224 397
rect 48 392 224 393
rect 275 403 276 407
rect 360 403 361 407
rect 275 402 361 403
rect 413 406 440 407
rect 413 402 414 406
rect 438 402 440 406
rect 275 397 396 402
rect 275 393 276 397
rect 395 393 396 397
rect 413 396 440 402
rect 413 392 414 396
rect 438 392 440 396
<< hvndcontact >>
rect 19 584 23 618
rect 39 614 173 618
rect 275 609 434 613
rect 39 604 173 608
rect 39 594 173 598
rect 39 584 173 588
rect 278 571 317 575
rect 15 546 19 570
rect 24 560 28 569
rect 24 551 28 555
rect 24 541 28 545
rect 33 541 37 570
rect 41 541 45 570
rect 50 560 54 564
rect 50 551 54 555
rect 50 541 54 545
rect 59 541 63 570
rect 68 560 72 564
rect 68 551 72 555
rect 68 541 72 545
rect 77 541 81 570
rect 86 560 90 564
rect 86 551 90 555
rect 86 541 90 545
rect 95 541 99 570
rect 104 560 108 564
rect 104 551 108 555
rect 104 541 108 545
rect 113 541 117 570
rect 122 560 126 564
rect 122 551 126 555
rect 122 541 126 545
rect 131 550 135 569
rect 140 541 144 570
rect 149 550 153 564
rect 149 541 153 545
rect 158 546 162 570
rect 167 541 171 570
rect 175 541 179 570
rect 184 560 188 569
rect 184 551 188 555
rect 184 541 188 545
rect 194 546 198 570
rect 202 541 206 570
rect 211 560 215 569
rect 211 551 215 555
rect 211 541 215 545
rect 221 546 225 570
rect 276 561 325 565
rect 276 551 325 555
rect 276 541 325 545
rect 330 541 334 570
rect 339 560 343 564
rect 339 551 343 555
rect 339 541 343 545
rect 348 541 352 570
rect 357 560 361 564
rect 357 551 361 555
rect 357 541 361 545
rect 366 541 370 570
rect 375 560 379 569
rect 375 551 379 555
rect 375 541 379 545
rect 384 541 388 570
rect 393 560 397 564
rect 393 551 397 555
rect 393 541 397 545
rect 402 541 406 570
rect 411 560 415 564
rect 411 551 415 555
rect 411 541 415 545
rect 420 541 424 570
rect 429 560 433 569
rect 429 551 433 555
rect 429 541 433 545
rect 50 352 174 356
rect 56 317 195 321
rect 56 311 195 315
rect 278 352 397 356
rect 51 276 185 280
rect 51 270 185 274
rect 255 317 394 321
rect 255 311 394 315
rect 265 276 399 280
rect 265 270 399 274
rect 56 230 195 239
rect 51 195 185 199
rect 51 189 185 193
rect 56 149 195 158
rect 255 230 394 239
rect 265 195 399 199
rect 265 189 399 193
rect 255 149 394 158
rect 51 114 185 118
rect 51 108 185 112
rect 56 68 195 77
rect 265 114 399 118
rect 265 108 399 112
rect 51 33 170 37
rect 255 68 394 77
rect 280 33 399 37
<< hvpdcontact >>
rect 41 972 170 976
rect 61 937 195 941
rect 61 931 195 935
rect 280 972 409 976
rect 255 937 389 941
rect 255 931 389 935
rect 46 896 190 900
rect 46 890 190 894
rect 260 896 404 900
rect 260 890 404 894
rect 61 850 195 859
rect 255 850 389 859
rect 46 815 190 819
rect 46 809 190 813
rect 61 769 195 778
rect 255 815 404 819
rect 260 809 404 813
rect 46 734 190 738
rect 46 728 190 732
rect 255 769 389 778
rect 260 734 404 738
rect 260 728 404 732
rect 61 688 195 697
rect 41 653 170 657
rect 255 688 389 697
rect 280 653 409 657
rect 276 473 325 477
rect 15 421 19 465
rect 24 462 28 466
rect 24 452 28 456
rect 24 442 28 446
rect 24 432 28 436
rect 33 422 37 471
rect 41 422 45 471
rect 50 462 54 466
rect 50 452 54 456
rect 50 442 54 446
rect 50 432 54 436
rect 59 422 63 471
rect 68 462 72 466
rect 68 452 72 456
rect 68 442 72 446
rect 68 432 72 436
rect 77 422 81 471
rect 86 462 90 466
rect 86 452 90 456
rect 86 442 90 446
rect 86 432 90 436
rect 95 422 99 471
rect 104 462 108 466
rect 104 452 108 456
rect 104 442 108 446
rect 104 432 108 436
rect 113 422 117 471
rect 122 462 126 466
rect 122 452 126 456
rect 122 442 126 446
rect 122 432 126 436
rect 131 422 135 471
rect 140 422 144 466
rect 149 466 153 470
rect 149 427 153 461
rect 158 422 162 471
rect 167 422 171 461
rect 176 422 180 471
rect 185 462 189 466
rect 185 452 189 456
rect 185 442 189 446
rect 185 432 189 436
rect 194 422 198 466
rect 203 422 207 471
rect 212 462 216 466
rect 212 452 216 456
rect 212 442 216 446
rect 212 432 216 436
rect 221 422 225 466
rect 276 463 325 467
rect 276 453 325 457
rect 276 443 325 447
rect 276 433 325 437
rect 276 423 325 427
rect 330 422 334 471
rect 339 462 343 466
rect 339 452 343 456
rect 339 441 343 445
rect 339 432 343 436
rect 348 427 352 471
rect 357 462 361 466
rect 357 452 361 456
rect 357 441 361 445
rect 357 432 361 436
rect 366 422 370 471
rect 375 462 379 466
rect 375 452 379 456
rect 375 441 379 445
rect 375 432 379 436
rect 384 422 388 471
rect 393 462 397 466
rect 393 452 397 456
rect 393 441 397 445
rect 393 432 397 436
rect 402 422 406 471
rect 411 466 415 470
rect 411 457 415 461
rect 411 447 415 451
rect 411 437 415 441
rect 411 427 415 431
rect 420 422 424 471
rect 276 413 325 417
rect 20 402 29 406
rect 429 408 433 472
rect 20 392 29 396
rect 49 393 223 397
rect 276 403 360 407
rect 414 402 438 406
rect 276 393 395 397
rect 414 392 438 396
<< hvpsubstratepdiff >>
rect 0 1008 450 1010
rect 0 1006 440 1008
rect 0 627 1 1006
rect 10 999 440 1006
rect 10 631 11 999
rect 439 631 440 999
rect 10 630 41 631
rect 10 627 14 630
rect 0 626 14 627
rect 28 627 41 630
rect 170 627 282 631
rect 436 629 440 631
rect 449 629 450 1008
rect 436 627 450 629
rect 28 626 450 627
rect 0 625 450 626
rect 0 521 6 625
rect 10 623 440 625
rect 10 619 275 623
rect 434 619 440 623
rect 10 618 440 619
rect 10 531 11 618
rect 437 603 440 618
rect 439 571 440 603
rect 50 531 54 533
rect 68 531 72 533
rect 86 531 90 533
rect 122 531 126 533
rect 275 531 325 533
rect 339 531 343 533
rect 357 531 361 533
rect 375 531 379 533
rect 393 531 397 533
rect 437 533 440 571
rect 411 531 415 533
rect 429 531 440 533
rect 10 530 440 531
rect 10 521 21 530
rect 25 526 41 530
rect 55 526 68 530
rect 92 526 105 530
rect 129 526 276 530
rect 345 526 356 530
rect 365 526 375 530
rect 399 526 409 530
rect 418 526 429 530
rect 438 526 440 530
rect 25 525 440 526
rect 25 521 188 525
rect 192 521 215 525
rect 219 521 440 525
rect 444 521 450 625
rect 0 520 450 521
rect 14 374 436 375
rect 14 365 20 374
rect 29 365 50 374
rect 14 360 50 365
rect 174 360 278 374
rect 397 365 421 374
rect 435 365 436 374
rect 397 360 436 365
rect 14 31 20 360
rect 24 359 426 360
rect 24 31 30 359
rect 38 357 213 359
rect 218 342 232 359
rect 237 357 412 359
rect 218 338 223 342
rect 227 338 232 342
rect 218 332 232 338
rect 218 323 223 332
rect 227 323 232 332
rect 218 317 232 323
rect 218 313 223 317
rect 227 313 232 317
rect 218 269 232 313
rect 218 265 223 269
rect 227 265 232 269
rect 218 259 232 265
rect 218 250 223 259
rect 227 250 232 259
rect 218 244 232 250
rect 218 235 223 244
rect 227 235 232 244
rect 218 229 232 235
rect 218 220 223 229
rect 227 220 232 229
rect 218 214 232 220
rect 218 210 223 214
rect 227 210 232 214
rect 218 172 232 210
rect 218 168 223 172
rect 227 168 232 172
rect 218 162 232 168
rect 218 153 223 162
rect 227 153 232 162
rect 218 147 232 153
rect 218 138 223 147
rect 227 138 232 147
rect 218 132 232 138
rect 218 123 223 132
rect 227 123 232 132
rect 218 117 232 123
rect 218 113 223 117
rect 227 113 232 117
rect 218 76 232 113
rect 218 72 223 76
rect 227 72 232 76
rect 218 66 232 72
rect 218 57 223 66
rect 227 57 232 66
rect 218 51 232 57
rect 218 47 223 51
rect 227 47 232 51
rect 14 30 30 31
rect 38 30 213 32
rect 218 30 232 47
rect 237 30 412 32
rect 420 31 426 359
rect 430 31 436 360
rect 14 26 416 30
rect 420 29 436 31
rect 14 22 50 26
rect 169 22 280 26
rect 399 25 416 26
rect 435 25 436 29
rect 399 22 436 25
rect 14 20 436 22
rect 14 16 20 20
rect 39 19 436 20
rect 39 16 421 19
rect 14 15 421 16
rect 435 15 436 19
rect 14 14 436 15
<< hvnsubstratendiff >>
rect 20 989 430 990
rect 24 988 430 989
rect 24 986 426 988
rect 24 982 280 986
rect 409 982 426 986
rect 24 981 426 982
rect 24 979 40 981
rect 24 650 30 979
rect 38 977 40 979
rect 174 979 426 981
rect 174 977 213 979
rect 218 925 232 979
rect 237 977 412 979
rect 218 921 223 925
rect 227 921 232 925
rect 218 915 232 921
rect 218 906 223 915
rect 227 906 232 915
rect 218 900 232 906
rect 218 891 223 900
rect 227 891 232 900
rect 218 885 232 891
rect 218 876 223 885
rect 227 876 232 885
rect 218 870 232 876
rect 218 866 223 870
rect 227 866 232 870
rect 218 834 232 866
rect 218 830 223 834
rect 227 830 232 834
rect 218 824 232 830
rect 218 815 223 824
rect 227 815 232 824
rect 218 809 232 815
rect 218 800 223 809
rect 227 800 232 809
rect 218 794 232 800
rect 218 785 223 794
rect 227 785 232 794
rect 218 779 232 785
rect 218 775 223 779
rect 227 775 232 779
rect 218 727 232 775
rect 218 723 223 727
rect 227 723 232 727
rect 218 717 232 723
rect 218 708 223 717
rect 227 708 232 717
rect 218 702 232 708
rect 218 693 223 702
rect 227 693 232 702
rect 218 687 232 693
rect 218 678 223 687
rect 227 678 232 687
rect 218 672 232 678
rect 218 668 223 672
rect 227 668 232 672
rect 38 651 213 652
rect 38 650 41 651
rect 24 645 41 650
rect 20 642 41 645
rect 140 650 213 651
rect 218 650 232 668
rect 237 651 412 652
rect 237 650 310 651
rect 140 642 310 650
rect 409 650 412 651
rect 420 650 426 979
rect 409 644 426 650
rect 409 642 430 644
rect 20 640 430 642
rect 0 489 450 490
rect 0 488 429 489
rect 0 484 2 488
rect 6 484 21 488
rect 25 484 46 488
rect 50 484 69 488
rect 73 484 79 488
rect 83 484 110 488
rect 114 484 120 488
rect 124 484 155 488
rect 159 484 188 488
rect 192 484 215 488
rect 219 487 429 488
rect 219 484 276 487
rect 0 483 276 484
rect 340 483 359 487
rect 363 483 375 487
rect 379 483 385 487
rect 389 483 395 487
rect 399 483 413 487
rect 417 485 429 487
rect 433 485 440 489
rect 417 483 440 485
rect 0 482 440 483
rect 0 479 8 482
rect 50 480 54 482
rect 68 480 72 482
rect 0 475 2 479
rect 6 475 8 479
rect 0 469 8 475
rect 86 480 90 482
rect 122 480 126 482
rect 275 478 325 482
rect 429 480 440 482
rect 0 465 2 469
rect 6 465 8 469
rect 0 459 8 465
rect 0 455 2 459
rect 6 455 8 459
rect 0 449 8 455
rect 0 445 2 449
rect 6 445 8 449
rect 0 439 8 445
rect 0 435 2 439
rect 6 435 8 439
rect 0 429 8 435
rect 0 425 2 429
rect 6 425 8 429
rect 0 419 8 425
rect 0 415 2 419
rect 6 415 8 419
rect 0 409 8 415
rect 0 405 2 409
rect 6 405 8 409
rect 0 399 8 405
rect 0 395 2 399
rect 6 395 8 399
rect 0 390 8 395
rect 13 390 30 392
rect 48 390 224 392
rect 275 390 396 393
rect 413 390 440 392
rect 0 389 440 390
rect 0 385 2 389
rect 6 386 440 389
rect 6 385 20 386
rect 0 382 20 385
rect 29 385 440 386
rect 444 385 450 489
rect 29 382 49 385
rect 0 381 49 382
rect 173 381 276 385
rect 395 381 414 385
rect 438 381 450 385
rect 0 2 2 381
rect 6 8 8 381
rect 442 8 444 381
rect 6 6 444 8
rect 6 2 10 6
rect 149 2 153 6
rect 297 2 301 6
rect 440 2 444 6
rect 448 2 450 381
rect 0 0 450 2
<< hvpsubstratepcontact >>
rect 1 627 10 1006
rect 14 626 28 630
rect 41 627 170 631
rect 282 627 436 631
rect 440 629 449 1008
rect 6 521 10 625
rect 275 619 434 623
rect 21 521 25 530
rect 41 526 55 530
rect 68 526 92 530
rect 105 526 129 530
rect 276 526 345 530
rect 356 526 365 530
rect 375 526 399 530
rect 409 526 418 530
rect 429 526 438 530
rect 188 521 192 525
rect 215 521 219 525
rect 440 521 444 625
rect 20 365 29 374
rect 50 360 174 374
rect 278 360 397 374
rect 421 365 435 374
rect 20 31 24 360
rect 223 338 227 342
rect 223 323 227 332
rect 223 313 227 317
rect 223 265 227 269
rect 223 250 227 259
rect 223 235 227 244
rect 223 220 227 229
rect 223 210 227 214
rect 223 168 227 172
rect 223 153 227 162
rect 223 138 227 147
rect 223 123 227 132
rect 223 113 227 117
rect 223 72 227 76
rect 223 57 227 66
rect 223 47 227 51
rect 426 31 430 360
rect 50 22 169 26
rect 280 22 399 26
rect 416 25 435 29
rect 20 16 39 20
rect 421 15 435 19
<< hvnsubstratencontact >>
rect 20 645 24 989
rect 280 982 409 986
rect 40 977 174 981
rect 223 921 227 925
rect 223 906 227 915
rect 223 891 227 900
rect 223 876 227 885
rect 223 866 227 870
rect 223 830 227 834
rect 223 815 227 824
rect 223 800 227 809
rect 223 785 227 794
rect 223 775 227 779
rect 223 723 227 727
rect 223 708 227 717
rect 223 693 227 702
rect 223 678 227 687
rect 223 668 227 672
rect 41 642 140 651
rect 310 642 409 651
rect 426 644 430 988
rect 2 484 6 488
rect 21 484 25 488
rect 46 484 50 488
rect 69 484 73 488
rect 79 484 83 488
rect 110 484 114 488
rect 120 484 124 488
rect 155 484 159 488
rect 188 484 192 488
rect 215 484 219 488
rect 276 483 340 487
rect 359 483 363 487
rect 375 483 379 487
rect 385 483 389 487
rect 395 483 399 487
rect 413 483 417 487
rect 429 485 433 489
rect 2 475 6 479
rect 2 465 6 469
rect 2 455 6 459
rect 2 445 6 449
rect 2 435 6 439
rect 2 425 6 429
rect 2 415 6 419
rect 2 405 6 409
rect 2 395 6 399
rect 2 385 6 389
rect 20 382 29 386
rect 440 385 444 489
rect 49 381 173 385
rect 276 381 395 385
rect 414 381 438 385
rect 2 2 6 381
rect 10 2 149 6
rect 153 2 297 6
rect 301 2 440 6
rect 444 2 448 381
<< polysilicon >>
rect 31 966 38 968
rect 31 742 32 966
rect 36 965 38 966
rect 213 965 216 968
rect 36 907 37 965
rect 234 965 237 968
rect 412 966 419 968
rect 412 965 414 966
rect 36 904 38 907
rect 213 904 216 907
rect 413 907 414 965
rect 36 886 37 904
rect 234 904 237 907
rect 412 904 414 907
rect 36 883 38 886
rect 213 883 216 886
rect 413 886 414 904
rect 36 826 37 883
rect 234 883 237 886
rect 412 883 414 886
rect 36 823 38 826
rect 213 823 216 826
rect 413 826 414 883
rect 36 805 37 823
rect 234 823 237 826
rect 412 823 414 826
rect 36 802 38 805
rect 213 802 216 805
rect 36 745 37 802
rect 413 805 414 823
rect 234 802 237 805
rect 412 802 414 805
rect 36 742 38 745
rect 213 742 216 745
rect 31 741 37 742
rect 413 745 414 802
rect 234 742 237 745
rect 412 742 414 745
rect 418 742 419 966
rect 31 723 38 724
rect 31 659 32 723
rect 36 721 38 723
rect 213 721 216 724
rect 413 741 419 742
rect 36 664 37 721
rect 234 721 237 724
rect 412 723 419 724
rect 412 721 414 723
rect 36 661 38 664
rect 213 661 216 664
rect 36 659 37 661
rect 31 658 37 659
rect 413 664 414 721
rect 234 661 237 664
rect 412 661 414 664
rect 413 659 414 661
rect 418 659 419 723
rect 413 658 419 659
rect 229 598 236 599
rect 229 594 230 598
rect 234 594 236 598
rect 229 592 236 594
rect 229 588 230 592
rect 234 588 236 592
rect 229 587 236 588
rect 429 598 436 599
rect 429 594 431 598
rect 435 594 436 598
rect 429 592 436 594
rect 429 588 431 592
rect 435 588 436 592
rect 429 587 436 588
rect 180 581 192 582
rect 19 580 30 581
rect 19 576 20 580
rect 29 576 30 580
rect 27 574 30 576
rect 180 577 182 581
rect 191 577 192 581
rect 180 576 192 577
rect 202 577 213 578
rect 20 570 23 573
rect 27 571 32 574
rect 29 570 32 571
rect 46 572 85 575
rect 46 570 49 572
rect 55 570 58 572
rect 64 570 67 572
rect 73 570 76 572
rect 82 570 85 572
rect 91 572 130 575
rect 91 570 94 572
rect 100 570 103 572
rect 109 570 112 572
rect 118 570 121 572
rect 127 570 130 572
rect 136 570 139 573
rect 145 570 148 573
rect 154 570 157 573
rect 163 570 166 573
rect 180 570 183 576
rect 202 573 203 577
rect 212 573 213 577
rect 371 577 377 578
rect 189 570 192 573
rect 202 572 213 573
rect 207 570 210 572
rect 216 570 219 573
rect 326 570 329 573
rect 335 572 347 575
rect 335 570 338 572
rect 344 570 347 572
rect 353 572 365 575
rect 353 570 356 572
rect 362 570 365 572
rect 371 573 372 577
rect 376 573 377 577
rect 371 572 377 573
rect 371 570 374 572
rect 380 570 383 573
rect 389 572 401 575
rect 389 570 392 572
rect 398 570 401 572
rect 407 572 419 575
rect 407 570 410 572
rect 416 570 419 572
rect 425 570 428 573
rect 20 539 23 540
rect 29 539 32 540
rect 13 538 23 539
rect 13 534 14 538
rect 18 536 23 538
rect 27 538 33 539
rect 18 534 19 536
rect 13 533 19 534
rect 27 534 28 538
rect 32 534 33 538
rect 46 537 49 540
rect 27 533 33 534
rect 55 539 58 540
rect 64 539 67 540
rect 55 538 67 539
rect 55 534 57 538
rect 66 534 67 538
rect 55 533 67 534
rect 73 537 76 540
rect 82 537 85 540
rect 91 539 94 540
rect 100 539 103 540
rect 91 538 103 539
rect 91 534 93 538
rect 102 534 103 538
rect 109 537 112 540
rect 118 537 121 540
rect 91 533 103 534
rect 127 537 130 540
rect 136 538 139 540
rect 145 538 148 540
rect 154 538 157 540
rect 163 538 166 540
rect 136 537 166 538
rect 136 535 151 537
rect 149 533 151 535
rect 160 535 166 537
rect 180 539 183 540
rect 189 539 192 540
rect 207 539 210 540
rect 216 539 219 540
rect 180 538 186 539
rect 160 533 161 535
rect 180 534 181 538
rect 185 534 186 538
rect 189 538 200 539
rect 189 536 195 538
rect 180 533 186 534
rect 194 534 195 536
rect 199 534 200 538
rect 194 533 200 534
rect 207 538 213 539
rect 207 534 208 538
rect 212 534 213 538
rect 216 538 227 539
rect 216 536 222 538
rect 207 533 213 534
rect 221 534 222 536
rect 226 534 227 538
rect 221 533 227 534
rect 326 539 329 540
rect 335 539 338 540
rect 326 536 338 539
rect 149 532 161 533
rect 344 539 347 540
rect 353 539 356 540
rect 344 536 356 539
rect 362 539 365 540
rect 371 539 374 540
rect 362 538 374 539
rect 362 534 363 538
rect 372 534 374 538
rect 362 533 374 534
rect 380 539 383 540
rect 389 539 392 540
rect 380 536 392 539
rect 398 539 401 540
rect 407 539 410 540
rect 398 536 410 539
rect 416 539 419 540
rect 425 539 428 540
rect 416 538 428 539
rect 416 534 418 538
rect 427 534 428 538
rect 416 533 428 534
rect 13 479 19 480
rect 13 475 14 479
rect 18 477 19 479
rect 27 479 33 480
rect 18 475 23 477
rect 13 474 23 475
rect 27 475 28 479
rect 32 475 33 479
rect 27 474 33 475
rect 20 472 23 474
rect 29 472 32 474
rect 46 472 49 475
rect 55 479 67 480
rect 55 475 57 479
rect 66 475 67 479
rect 55 474 67 475
rect 55 472 58 474
rect 64 472 67 474
rect 73 472 76 475
rect 82 472 85 475
rect 91 479 103 480
rect 91 475 92 479
rect 101 475 103 479
rect 91 474 103 475
rect 91 472 94 474
rect 100 472 103 474
rect 109 472 112 475
rect 118 472 121 475
rect 140 480 151 481
rect 140 477 141 480
rect 136 476 141 477
rect 150 477 151 480
rect 180 479 186 480
rect 150 476 166 477
rect 127 472 130 475
rect 136 474 166 476
rect 180 475 181 479
rect 185 475 186 479
rect 194 479 200 480
rect 194 477 195 479
rect 180 474 186 475
rect 190 475 195 477
rect 199 475 200 479
rect 190 474 200 475
rect 207 479 213 480
rect 207 475 208 479
rect 212 475 213 479
rect 221 479 227 480
rect 221 477 222 479
rect 207 474 213 475
rect 217 475 222 477
rect 226 475 227 479
rect 217 474 227 475
rect 362 479 374 480
rect 136 472 139 474
rect 145 472 148 474
rect 154 472 157 474
rect 163 472 166 474
rect 181 472 184 474
rect 190 472 193 474
rect 208 472 211 474
rect 217 472 220 474
rect 326 474 338 477
rect 326 472 329 474
rect 335 472 338 474
rect 344 474 356 477
rect 344 472 347 474
rect 353 472 356 474
rect 362 475 364 479
rect 373 475 374 479
rect 416 479 428 480
rect 362 474 374 475
rect 362 472 365 474
rect 371 472 374 474
rect 380 474 392 477
rect 380 472 383 474
rect 389 472 392 474
rect 398 474 410 477
rect 398 472 401 474
rect 407 472 410 474
rect 416 475 418 479
rect 427 475 428 479
rect 416 474 428 475
rect 416 472 419 474
rect 425 472 428 474
rect 20 419 23 420
rect 29 419 32 420
rect 46 419 49 420
rect 55 419 58 420
rect 12 418 23 419
rect 12 414 13 418
rect 22 414 23 418
rect 12 413 23 414
rect 26 418 37 419
rect 26 414 27 418
rect 36 414 37 418
rect 26 413 37 414
rect 46 418 58 419
rect 46 414 47 418
rect 56 415 58 418
rect 64 415 67 420
rect 73 415 76 420
rect 82 415 85 420
rect 56 414 85 415
rect 46 412 85 414
rect 91 415 94 420
rect 100 415 103 420
rect 109 415 112 420
rect 118 415 121 420
rect 127 415 130 420
rect 136 417 139 420
rect 145 417 148 420
rect 154 417 157 420
rect 163 417 166 420
rect 181 419 184 420
rect 176 418 187 419
rect 91 412 130 415
rect 176 414 177 418
rect 186 414 187 418
rect 190 417 193 420
rect 208 415 211 420
rect 217 417 220 420
rect 326 417 329 420
rect 335 419 338 420
rect 344 419 347 420
rect 176 413 187 414
rect 206 414 211 415
rect 206 410 207 414
rect 216 410 217 414
rect 206 409 217 410
rect 335 416 347 419
rect 353 419 356 420
rect 362 419 365 420
rect 353 416 365 419
rect 371 417 374 420
rect 380 417 383 420
rect 389 419 392 420
rect 398 419 401 420
rect 389 416 401 419
rect 407 419 410 420
rect 416 419 419 420
rect 407 416 419 419
rect 425 417 428 420
rect 31 348 37 349
rect 31 344 32 348
rect 36 345 38 348
rect 213 345 216 348
rect 36 344 37 345
rect 31 343 37 344
rect 413 349 419 350
rect 413 348 414 349
rect 234 345 237 348
rect 412 345 414 348
rect 418 345 419 349
rect 31 286 38 287
rect 31 42 32 286
rect 36 284 38 286
rect 213 284 216 287
rect 36 266 37 284
rect 413 344 419 345
rect 234 284 237 287
rect 412 286 419 287
rect 412 284 414 286
rect 36 263 38 266
rect 213 263 216 266
rect 413 266 414 284
rect 36 206 37 263
rect 234 263 237 266
rect 412 263 414 266
rect 36 203 38 206
rect 213 203 216 206
rect 36 185 37 203
rect 36 182 38 185
rect 213 182 216 185
rect 36 125 37 182
rect 413 206 414 263
rect 234 203 237 206
rect 412 203 414 206
rect 413 185 414 203
rect 234 182 237 185
rect 412 182 414 185
rect 36 122 38 125
rect 213 122 216 125
rect 413 125 414 182
rect 36 104 37 122
rect 234 122 237 125
rect 412 122 414 125
rect 36 101 38 104
rect 213 101 216 104
rect 36 44 37 101
rect 413 104 414 122
rect 234 101 237 104
rect 412 101 414 104
rect 36 42 38 44
rect 31 41 38 42
rect 213 41 216 44
rect 413 44 414 101
rect 234 41 237 44
rect 412 42 414 44
rect 418 42 419 286
rect 412 41 419 42
<< polycontact >>
rect 32 742 36 966
rect 414 742 418 966
rect 32 659 36 723
rect 414 659 418 723
rect 230 594 234 598
rect 230 588 234 592
rect 431 594 435 598
rect 431 588 435 592
rect 20 576 29 580
rect 182 577 191 581
rect 203 573 212 577
rect 372 573 376 577
rect 14 534 18 538
rect 28 534 32 538
rect 57 534 66 538
rect 93 534 102 538
rect 151 533 160 537
rect 181 534 185 538
rect 195 534 199 538
rect 208 534 212 538
rect 222 534 226 538
rect 363 534 372 538
rect 418 534 427 538
rect 14 475 18 479
rect 28 475 32 479
rect 57 475 66 479
rect 92 475 101 479
rect 141 476 150 480
rect 181 475 185 479
rect 195 475 199 479
rect 208 475 212 479
rect 222 475 226 479
rect 364 475 373 479
rect 418 475 427 479
rect 13 414 22 418
rect 27 414 36 418
rect 47 414 56 418
rect 177 414 186 418
rect 207 410 216 414
rect 32 344 36 348
rect 414 345 418 349
rect 32 42 36 286
rect 414 42 418 286
<< metal1 >>
rect 30 1495 420 1500
rect 30 1114 34 1495
rect 415 1114 420 1495
rect 30 1110 420 1114
rect 137 1100 313 1110
rect 147 1090 303 1100
rect 157 1080 293 1090
rect 167 1070 283 1080
rect 0 1006 174 1010
rect 0 627 1 1006
rect 10 999 174 1006
rect 10 631 11 999
rect 178 998 272 1070
rect 276 1008 450 1010
rect 276 999 440 1008
rect 24 988 173 989
rect 24 987 174 988
rect 24 648 25 987
rect 29 986 174 987
rect 29 982 40 986
rect 181 984 269 998
rect 277 988 430 989
rect 276 987 426 988
rect 276 986 421 987
rect 29 981 174 982
rect 29 977 40 981
rect 29 976 174 977
rect 29 972 41 976
rect 170 972 174 976
rect 29 966 174 972
rect 186 969 264 984
rect 276 982 280 986
rect 409 982 421 986
rect 276 981 421 982
rect 276 977 280 981
rect 409 977 421 981
rect 276 976 421 977
rect 276 972 280 976
rect 409 972 421 976
rect 29 742 32 966
rect 36 964 174 966
rect 36 940 39 964
rect 48 960 52 964
rect 171 960 174 964
rect 48 940 51 960
rect 199 957 251 969
rect 276 966 421 972
rect 276 964 414 966
rect 276 960 284 964
rect 398 960 402 964
rect 36 932 51 940
rect 36 908 39 932
rect 48 912 51 932
rect 56 941 394 957
rect 56 937 61 941
rect 195 937 255 941
rect 389 937 394 941
rect 56 935 394 937
rect 56 931 61 935
rect 195 931 255 935
rect 389 931 394 935
rect 56 928 394 931
rect 56 915 220 928
rect 48 908 52 912
rect 191 908 195 912
rect 36 900 195 908
rect 36 896 46 900
rect 190 896 195 900
rect 36 894 195 896
rect 36 890 46 894
rect 190 890 195 894
rect 36 882 195 890
rect 36 858 39 882
rect 48 878 52 882
rect 191 878 195 882
rect 48 858 51 878
rect 199 875 220 915
rect 36 851 51 858
rect 36 827 39 851
rect 48 831 51 851
rect 56 863 220 875
rect 223 920 227 921
rect 223 915 227 916
rect 223 905 227 906
rect 223 900 227 901
rect 223 890 227 891
rect 223 885 227 886
rect 223 875 227 876
rect 223 870 227 871
rect 230 915 394 928
rect 399 940 402 960
rect 411 940 414 964
rect 399 932 414 940
rect 230 875 251 915
rect 399 912 402 932
rect 255 908 264 912
rect 398 908 402 912
rect 411 908 414 932
rect 255 900 414 908
rect 255 896 260 900
rect 404 896 414 900
rect 255 894 414 896
rect 255 890 260 894
rect 404 890 414 894
rect 255 882 414 890
rect 255 878 264 882
rect 398 878 402 882
rect 230 863 394 875
rect 56 859 394 863
rect 56 850 61 859
rect 195 850 255 859
rect 389 850 394 859
rect 56 837 394 850
rect 56 834 220 837
rect 230 834 394 837
rect 399 858 402 878
rect 411 858 414 882
rect 399 851 414 858
rect 48 827 52 831
rect 191 827 195 831
rect 36 819 195 827
rect 36 815 46 819
rect 190 815 195 819
rect 36 813 195 815
rect 36 809 46 813
rect 190 809 195 813
rect 36 801 195 809
rect 36 777 39 801
rect 48 797 52 801
rect 191 797 195 801
rect 48 777 51 797
rect 199 794 220 834
rect 36 770 51 777
rect 36 746 39 770
rect 48 750 51 770
rect 56 778 220 794
rect 56 769 61 778
rect 195 772 220 778
rect 223 829 227 830
rect 223 824 227 825
rect 223 814 227 815
rect 223 809 227 810
rect 223 799 227 800
rect 223 794 227 795
rect 223 784 227 785
rect 223 779 227 780
rect 230 794 251 834
rect 399 831 402 851
rect 255 827 259 831
rect 398 827 402 831
rect 411 827 414 851
rect 255 819 414 827
rect 404 815 414 819
rect 255 813 414 815
rect 255 809 260 813
rect 404 809 414 813
rect 255 801 414 809
rect 255 797 259 801
rect 398 797 402 801
rect 230 778 394 794
rect 230 772 255 778
rect 195 769 255 772
rect 389 769 394 778
rect 56 753 394 769
rect 399 777 402 797
rect 411 777 414 801
rect 399 770 414 777
rect 48 746 52 750
rect 191 746 195 750
rect 36 742 195 746
rect 39 738 195 742
rect 39 734 46 738
rect 190 734 195 738
rect 39 732 195 734
rect 39 728 46 732
rect 190 728 195 732
rect 24 645 29 648
rect 20 641 29 645
rect 32 723 36 724
rect 32 645 36 659
rect 39 720 195 728
rect 48 716 52 720
rect 191 716 195 720
rect 199 730 251 753
rect 399 750 402 770
rect 48 696 51 716
rect 199 713 220 730
rect 39 689 51 696
rect 48 669 51 689
rect 56 697 220 713
rect 56 688 61 697
rect 195 688 220 697
rect 56 672 220 688
rect 48 665 52 669
rect 171 665 174 669
rect 39 657 174 665
rect 39 653 41 657
rect 170 653 174 657
rect 39 651 174 653
rect 39 642 41 651
rect 140 642 174 651
rect 39 641 174 642
rect 178 665 220 672
rect 223 722 227 723
rect 223 717 227 718
rect 223 707 227 708
rect 223 702 227 703
rect 223 692 227 693
rect 223 687 227 688
rect 223 677 227 678
rect 223 672 227 673
rect 230 713 251 730
rect 255 746 259 750
rect 398 746 402 750
rect 411 746 414 770
rect 255 742 414 746
rect 418 742 421 966
rect 255 738 411 742
rect 255 734 260 738
rect 404 734 411 738
rect 255 732 411 734
rect 255 728 260 732
rect 404 728 411 732
rect 255 720 411 728
rect 255 716 259 720
rect 398 716 402 720
rect 230 697 394 713
rect 230 688 255 697
rect 389 688 394 697
rect 230 672 394 688
rect 399 696 402 716
rect 399 689 411 696
rect 230 665 272 672
rect 399 669 402 689
rect 32 636 36 641
rect 10 630 29 631
rect 10 627 14 630
rect 0 626 14 627
rect 28 626 29 630
rect 0 625 29 626
rect 0 521 1 625
rect 5 521 6 625
rect 10 621 14 625
rect 28 621 29 625
rect 10 618 29 621
rect 10 584 14 618
rect 18 584 19 618
rect 23 584 24 618
rect 28 584 29 618
rect 10 521 11 584
rect 32 580 36 632
rect 39 627 41 630
rect 170 627 174 631
rect 39 623 174 627
rect 173 620 174 623
rect 39 618 173 619
rect 39 613 173 614
rect 39 608 173 609
rect 39 603 173 604
rect 39 598 173 599
rect 39 593 173 594
rect 39 588 173 589
rect 178 598 272 665
rect 276 665 279 669
rect 398 665 402 669
rect 276 657 411 665
rect 276 653 280 657
rect 409 653 411 657
rect 276 651 411 653
rect 276 642 310 651
rect 409 642 411 651
rect 276 641 411 642
rect 414 645 418 659
rect 425 648 426 987
rect 421 644 426 648
rect 414 638 418 641
rect 439 631 440 999
rect 276 627 282 631
rect 436 629 440 631
rect 449 629 450 1008
rect 436 627 450 629
rect 276 625 450 627
rect 276 624 440 625
rect 275 623 440 624
rect 434 619 440 623
rect 275 618 440 619
rect 434 614 440 618
rect 275 613 440 614
rect 434 609 440 613
rect 275 608 440 609
rect 434 604 440 608
rect 437 603 440 604
rect 178 594 230 598
rect 234 594 272 598
rect 178 592 272 594
rect 178 588 230 592
rect 234 588 272 592
rect 178 586 272 588
rect 431 592 435 594
rect 431 587 435 588
rect 16 576 20 579
rect 32 576 179 580
rect 191 577 198 580
rect 16 570 19 576
rect 41 570 135 572
rect 24 569 28 570
rect 24 555 28 556
rect 24 550 28 551
rect 24 545 28 546
rect 22 541 24 544
rect 37 541 38 546
rect 45 568 59 570
rect 50 564 54 565
rect 50 555 54 556
rect 50 550 54 551
rect 50 545 54 546
rect 63 568 77 570
rect 68 564 72 565
rect 68 555 72 556
rect 68 550 72 551
rect 68 545 72 546
rect 81 568 95 570
rect 86 564 90 565
rect 86 555 90 556
rect 86 550 90 551
rect 86 545 90 546
rect 99 568 113 570
rect 104 564 108 565
rect 104 555 108 556
rect 104 550 108 551
rect 104 545 108 546
rect 117 569 135 570
rect 117 568 131 569
rect 122 564 126 565
rect 122 555 126 556
rect 122 550 126 551
rect 140 570 162 572
rect 175 570 179 576
rect 194 570 198 577
rect 212 573 225 577
rect 221 570 225 573
rect 122 545 126 546
rect 0 488 7 489
rect 0 480 2 488
rect 6 480 7 488
rect 0 479 7 480
rect 0 475 2 479
rect 6 475 7 479
rect 14 479 18 534
rect 22 530 25 541
rect 28 512 32 534
rect 0 474 7 475
rect 0 470 2 474
rect 6 470 7 474
rect 0 469 7 470
rect 0 465 2 469
rect 6 465 7 469
rect 22 471 25 484
rect 28 479 32 503
rect 35 499 38 541
rect 50 538 54 541
rect 69 538 72 541
rect 86 538 90 541
rect 122 538 126 541
rect 132 541 140 543
rect 144 568 158 570
rect 132 539 144 541
rect 149 564 153 565
rect 149 545 153 546
rect 153 541 167 543
rect 149 540 171 541
rect 41 531 54 538
rect 41 530 55 531
rect 41 525 55 526
rect 35 471 38 495
rect 45 484 46 488
rect 50 484 51 488
rect 41 482 55 484
rect 41 474 54 482
rect 58 479 61 534
rect 69 531 90 538
rect 69 530 92 531
rect 68 525 92 526
rect 95 507 99 534
rect 105 530 129 538
rect 105 525 129 526
rect 132 515 135 539
rect 68 484 69 488
rect 73 484 74 488
rect 78 484 79 488
rect 83 484 84 488
rect 88 484 89 488
rect 64 483 89 484
rect 50 471 54 474
rect 69 474 89 483
rect 92 479 101 495
rect 104 484 105 488
rect 109 484 110 488
rect 114 484 115 488
rect 119 484 120 488
rect 124 484 125 488
rect 104 475 129 484
rect 69 471 72 474
rect 86 471 89 474
rect 122 471 126 475
rect 132 472 135 511
rect 143 480 147 503
rect 155 499 159 533
rect 167 503 171 540
rect 154 484 155 488
rect 159 484 160 488
rect 167 472 171 494
rect 132 471 153 472
rect 22 467 24 471
rect 24 466 28 467
rect 0 464 7 465
rect 0 460 2 464
rect 6 460 7 464
rect 0 459 7 460
rect 0 455 2 459
rect 6 455 7 459
rect 0 454 7 455
rect 0 450 2 454
rect 6 450 7 454
rect 0 449 7 450
rect 0 445 2 449
rect 6 445 7 449
rect 0 444 7 445
rect 0 440 2 444
rect 6 440 7 444
rect 0 439 7 440
rect 0 435 2 439
rect 6 435 7 439
rect 0 434 7 435
rect 0 430 2 434
rect 6 430 7 434
rect 0 429 7 430
rect 0 425 2 429
rect 6 425 7 429
rect 0 424 7 425
rect 0 420 2 424
rect 6 420 7 424
rect 24 461 28 462
rect 24 456 28 457
rect 24 451 28 452
rect 24 446 28 447
rect 24 441 28 442
rect 24 436 28 437
rect 24 431 28 432
rect 19 421 29 424
rect 37 463 38 471
rect 50 466 54 467
rect 50 461 54 462
rect 50 456 54 457
rect 50 451 54 452
rect 50 446 54 447
rect 50 441 54 442
rect 50 436 54 437
rect 50 431 54 432
rect 45 422 59 424
rect 68 466 72 467
rect 68 461 72 462
rect 68 456 72 457
rect 68 451 72 452
rect 68 446 72 447
rect 68 441 72 442
rect 68 436 72 437
rect 68 431 72 432
rect 41 421 63 422
rect 0 419 7 420
rect 0 415 2 419
rect 6 415 7 419
rect 25 418 29 421
rect 59 420 63 421
rect 86 466 90 467
rect 86 461 90 462
rect 86 456 90 457
rect 86 451 90 452
rect 86 446 90 447
rect 86 441 90 442
rect 86 436 90 437
rect 86 431 90 432
rect 77 420 81 422
rect 104 466 108 467
rect 104 461 108 462
rect 104 456 108 457
rect 104 451 108 452
rect 104 446 108 447
rect 104 441 108 442
rect 104 436 108 437
rect 104 431 108 432
rect 95 420 99 422
rect 122 466 126 467
rect 122 461 126 462
rect 122 456 126 457
rect 122 451 126 452
rect 122 446 126 447
rect 122 441 126 442
rect 122 436 126 437
rect 122 431 126 432
rect 113 420 117 422
rect 135 470 153 471
rect 135 469 149 470
rect 131 420 135 422
rect 149 461 153 462
rect 158 471 171 472
rect 144 422 158 424
rect 162 469 171 471
rect 184 569 188 570
rect 184 555 188 556
rect 184 550 188 551
rect 184 545 188 546
rect 175 471 178 541
rect 181 479 185 534
rect 188 530 191 544
rect 211 569 215 570
rect 211 555 215 556
rect 211 550 215 551
rect 211 545 215 546
rect 188 525 192 526
rect 195 515 199 534
rect 188 471 191 484
rect 195 479 199 511
rect 175 463 176 471
rect 167 461 171 462
rect 189 468 191 471
rect 202 471 205 541
rect 208 479 212 534
rect 215 530 218 544
rect 215 525 219 526
rect 222 503 226 534
rect 215 471 218 484
rect 222 479 226 494
rect 185 466 189 467
rect 185 461 189 462
rect 185 456 189 457
rect 185 451 189 452
rect 185 446 189 447
rect 185 441 189 442
rect 185 436 189 437
rect 185 431 189 432
rect 184 422 194 424
rect 202 463 203 471
rect 140 421 162 422
rect 0 414 7 415
rect 0 410 2 414
rect 6 410 7 414
rect 0 409 7 410
rect 0 405 2 409
rect 6 405 7 409
rect 0 404 7 405
rect 0 400 2 404
rect 6 400 7 404
rect 0 399 7 400
rect 0 395 2 399
rect 6 395 7 399
rect 0 394 7 395
rect 0 390 2 394
rect 6 390 7 394
rect 0 389 7 390
rect 25 414 27 418
rect 42 414 47 418
rect 59 416 135 420
rect 184 420 198 422
rect 201 422 203 430
rect 216 468 218 471
rect 212 466 216 467
rect 212 461 216 462
rect 212 456 216 457
rect 212 451 216 452
rect 212 446 216 447
rect 212 441 216 442
rect 212 436 216 437
rect 212 431 216 432
rect 212 422 221 424
rect 184 418 187 420
rect 186 414 187 418
rect 201 417 204 422
rect 0 385 2 389
rect 6 385 8 389
rect 0 381 8 385
rect 0 2 2 381
rect 6 6 8 381
rect 13 13 17 414
rect 20 406 29 407
rect 20 401 29 402
rect 20 396 29 397
rect 20 391 29 392
rect 20 386 29 387
rect 20 381 29 382
rect 20 374 29 375
rect 20 360 29 365
rect 24 31 25 360
rect 32 374 36 407
rect 32 348 36 365
rect 29 42 32 286
rect 36 42 38 286
rect 29 31 38 42
rect 20 25 38 31
rect 20 20 39 21
rect 42 13 46 414
rect 190 413 204 417
rect 212 420 225 422
rect 212 414 216 420
rect 190 411 194 413
rect 53 407 194 411
rect 49 402 223 404
rect 49 397 223 398
rect 49 391 223 393
rect 49 385 173 387
rect 229 386 272 586
rect 372 582 435 587
rect 276 580 320 581
rect 276 576 278 580
rect 317 576 320 580
rect 276 575 320 576
rect 276 571 278 575
rect 317 571 320 575
rect 330 576 369 580
rect 276 570 325 571
rect 276 565 325 566
rect 276 560 325 561
rect 276 555 325 556
rect 276 550 325 551
rect 276 545 325 546
rect 330 570 334 576
rect 348 570 352 576
rect 339 564 343 565
rect 339 555 343 556
rect 339 550 343 551
rect 339 545 343 546
rect 276 540 325 541
rect 276 535 325 536
rect 339 535 343 541
rect 366 570 369 576
rect 372 577 377 582
rect 376 573 377 577
rect 384 576 424 579
rect 384 570 388 576
rect 276 530 345 535
rect 276 525 345 526
rect 348 510 352 541
rect 357 564 361 565
rect 357 555 361 556
rect 357 550 361 551
rect 357 545 361 546
rect 375 569 379 570
rect 375 555 379 556
rect 375 550 379 551
rect 375 545 379 546
rect 402 570 406 576
rect 393 564 397 565
rect 393 555 397 556
rect 393 550 397 551
rect 393 545 397 546
rect 357 531 360 541
rect 355 530 365 531
rect 355 526 356 530
rect 355 525 365 526
rect 355 521 356 525
rect 275 483 276 487
rect 340 483 343 487
rect 275 482 325 483
rect 275 478 276 482
rect 275 477 325 478
rect 275 473 276 477
rect 275 472 325 473
rect 275 468 276 472
rect 339 471 343 483
rect 275 467 325 468
rect 275 463 276 467
rect 275 462 325 463
rect 275 458 276 462
rect 275 457 325 458
rect 275 453 276 457
rect 275 452 325 453
rect 275 448 276 452
rect 275 447 325 448
rect 275 443 276 447
rect 275 442 325 443
rect 275 438 276 442
rect 275 437 325 438
rect 275 433 276 437
rect 275 432 325 433
rect 275 428 276 432
rect 49 374 174 375
rect 49 360 50 374
rect 49 356 174 360
rect 49 352 50 356
rect 49 344 174 352
rect 53 340 57 344
rect 171 340 174 344
rect 178 345 272 386
rect 276 427 325 428
rect 276 422 325 423
rect 276 417 325 418
rect 276 412 325 413
rect 339 466 343 467
rect 339 461 343 462
rect 339 456 343 457
rect 339 451 343 452
rect 339 445 343 447
rect 339 436 343 437
rect 339 431 343 432
rect 348 471 352 501
rect 357 471 361 483
rect 368 479 372 534
rect 375 535 379 541
rect 393 535 397 541
rect 420 570 424 576
rect 439 571 440 603
rect 437 570 440 571
rect 375 530 399 535
rect 375 525 399 526
rect 379 483 380 487
rect 384 483 385 487
rect 389 483 390 487
rect 394 483 395 487
rect 376 471 379 483
rect 393 471 397 483
rect 357 466 361 467
rect 357 461 361 462
rect 357 456 361 457
rect 357 451 361 452
rect 357 445 361 447
rect 357 436 361 437
rect 357 431 361 432
rect 330 414 334 422
rect 348 414 352 427
rect 375 466 379 467
rect 375 461 379 462
rect 375 456 379 457
rect 375 451 379 452
rect 375 445 379 447
rect 375 436 379 437
rect 375 431 379 432
rect 393 466 397 467
rect 393 461 397 462
rect 393 456 397 457
rect 393 451 397 452
rect 393 445 397 447
rect 393 436 397 437
rect 393 431 397 432
rect 402 471 406 541
rect 411 564 415 565
rect 411 555 415 556
rect 411 550 415 551
rect 411 545 415 546
rect 429 569 440 570
rect 433 556 440 569
rect 429 555 440 556
rect 433 551 440 555
rect 429 550 440 551
rect 433 546 440 550
rect 429 545 440 546
rect 433 541 440 545
rect 411 531 415 541
rect 409 530 418 531
rect 409 525 418 526
rect 421 510 425 534
rect 430 531 440 541
rect 429 530 440 531
rect 438 526 440 530
rect 429 525 440 526
rect 438 521 440 525
rect 444 521 445 625
rect 449 521 450 625
rect 366 414 370 422
rect 330 411 370 414
rect 384 415 388 422
rect 411 470 415 483
rect 421 479 425 501
rect 433 485 434 489
rect 438 485 440 489
rect 430 477 440 485
rect 430 472 434 477
rect 411 461 415 462
rect 411 456 415 457
rect 411 451 415 452
rect 411 446 415 447
rect 411 441 415 442
rect 411 436 415 437
rect 411 431 415 432
rect 402 415 406 422
rect 420 415 424 422
rect 384 411 424 415
rect 366 408 370 411
rect 276 407 360 408
rect 366 404 405 408
rect 276 402 360 403
rect 360 398 395 401
rect 276 397 395 398
rect 276 391 395 393
rect 276 385 395 387
rect 178 337 220 345
rect 49 312 53 320
rect 56 321 220 337
rect 195 317 220 321
rect 56 315 220 317
rect 195 311 220 315
rect 223 337 227 338
rect 223 332 227 333
rect 223 322 227 323
rect 223 317 227 318
rect 230 337 272 345
rect 276 374 399 375
rect 276 360 278 374
rect 397 360 399 374
rect 276 356 399 360
rect 276 352 278 356
rect 397 352 399 356
rect 276 344 399 352
rect 276 340 277 344
rect 396 340 399 344
rect 230 321 394 337
rect 230 317 255 321
rect 230 315 394 317
rect 56 310 220 311
rect 230 311 255 315
rect 230 310 394 311
rect 56 295 394 310
rect 53 288 57 292
rect 181 288 185 292
rect 49 280 185 288
rect 49 276 51 280
rect 49 274 185 276
rect 49 270 51 274
rect 49 262 185 270
rect 53 258 57 262
rect 181 258 185 262
rect 189 272 261 295
rect 189 255 220 272
rect 49 231 53 238
rect 56 239 220 255
rect 195 230 220 239
rect 56 214 220 230
rect 53 207 57 211
rect 181 207 185 211
rect 49 199 185 207
rect 49 195 51 199
rect 49 193 185 195
rect 49 189 51 193
rect 49 181 185 189
rect 53 177 57 181
rect 181 177 185 181
rect 189 207 220 214
rect 223 264 227 265
rect 223 259 227 260
rect 223 249 227 250
rect 223 244 227 245
rect 223 234 227 235
rect 223 229 227 230
rect 223 219 227 220
rect 223 214 227 215
rect 230 255 261 272
rect 265 288 267 292
rect 396 288 399 292
rect 265 280 399 288
rect 265 274 399 276
rect 265 262 399 270
rect 265 258 267 262
rect 396 258 399 262
rect 230 239 394 255
rect 230 230 255 239
rect 230 214 394 230
rect 230 207 261 214
rect 189 175 261 207
rect 265 207 267 211
rect 396 207 399 211
rect 265 199 399 207
rect 265 193 399 195
rect 265 181 399 189
rect 265 177 267 181
rect 396 177 399 181
rect 189 174 220 175
rect 49 150 53 157
rect 56 158 220 174
rect 230 174 261 175
rect 195 149 220 158
rect 56 133 220 149
rect 53 126 57 130
rect 181 126 185 130
rect 49 118 185 126
rect 49 114 51 118
rect 49 112 185 114
rect 49 108 51 112
rect 49 100 185 108
rect 53 96 57 100
rect 181 96 185 100
rect 189 110 220 133
rect 223 167 227 168
rect 223 162 227 163
rect 223 152 227 153
rect 223 147 227 148
rect 223 137 227 138
rect 223 132 227 133
rect 223 122 227 123
rect 223 117 227 118
rect 230 158 394 174
rect 230 149 255 158
rect 230 133 394 149
rect 230 110 261 133
rect 189 93 261 110
rect 265 126 267 130
rect 396 126 399 130
rect 265 118 399 126
rect 265 112 399 114
rect 265 100 399 108
rect 265 96 267 100
rect 396 96 399 100
rect 49 69 53 76
rect 56 79 394 93
rect 56 77 220 79
rect 195 68 220 77
rect 230 77 394 79
rect 56 52 220 68
rect 53 45 57 49
rect 171 45 174 49
rect 49 37 174 45
rect 49 33 51 37
rect 170 33 174 37
rect 49 31 174 33
rect 49 27 50 31
rect 169 27 174 31
rect 49 26 174 27
rect 49 22 50 26
rect 169 22 174 26
rect 49 21 174 22
rect 49 17 50 21
rect 169 17 174 21
rect 49 16 174 17
rect 63 14 174 16
rect 177 44 220 52
rect 223 71 227 72
rect 223 66 227 67
rect 223 56 227 57
rect 223 51 227 52
rect 230 68 255 77
rect 230 52 394 68
rect 230 44 273 52
rect 177 29 273 44
rect 177 15 178 29
rect 272 15 273 29
rect 177 14 273 15
rect 276 45 277 49
rect 396 45 399 49
rect 276 37 399 45
rect 276 33 280 37
rect 276 31 399 33
rect 276 27 280 31
rect 276 26 399 27
rect 276 22 280 26
rect 276 21 399 22
rect 276 17 280 21
rect 276 16 399 17
rect 276 14 392 16
rect 402 13 405 404
rect 404 9 405 13
rect 408 13 411 411
rect 433 408 434 472
rect 438 408 440 477
rect 429 407 440 408
rect 414 406 440 407
rect 438 402 440 406
rect 414 401 440 402
rect 438 397 440 401
rect 414 396 440 397
rect 438 392 440 396
rect 414 391 440 392
rect 438 387 440 391
rect 414 385 440 387
rect 444 385 445 489
rect 449 385 450 489
rect 438 381 450 385
rect 421 374 436 375
rect 414 349 418 365
rect 435 365 436 374
rect 421 360 436 365
rect 418 42 421 286
rect 414 31 421 42
rect 425 31 426 360
rect 430 31 431 360
rect 435 31 436 360
rect 414 29 436 31
rect 414 25 416 29
rect 435 25 436 29
rect 414 24 436 25
rect 414 20 416 24
rect 435 20 436 24
rect 414 19 436 20
rect 414 16 421 19
rect 420 15 421 16
rect 435 15 436 19
rect 420 14 436 15
rect 442 8 444 381
rect 23 6 35 8
rect 51 6 392 8
rect 420 6 444 8
rect 6 2 10 6
rect 149 2 153 6
rect 297 2 301 6
rect 440 2 444 6
rect 448 2 450 381
rect 0 0 450 2
<< m2contact >>
rect 25 648 29 987
rect 40 982 174 986
rect 280 977 409 981
rect 39 940 48 964
rect 52 960 171 964
rect 284 960 398 964
rect 39 908 48 932
rect 52 908 191 912
rect 39 858 48 882
rect 52 878 191 882
rect 39 827 48 851
rect 223 916 227 920
rect 223 901 227 905
rect 223 886 227 890
rect 223 871 227 875
rect 402 940 411 964
rect 264 908 398 912
rect 402 908 411 932
rect 264 878 398 882
rect 402 858 411 882
rect 52 827 191 831
rect 39 777 48 801
rect 52 797 191 801
rect 39 746 48 770
rect 223 825 227 829
rect 223 810 227 814
rect 223 795 227 799
rect 223 780 227 784
rect 259 827 398 831
rect 402 827 411 851
rect 259 797 398 801
rect 402 777 411 801
rect 52 746 191 750
rect 32 641 36 645
rect 39 696 48 720
rect 52 716 191 720
rect 39 665 48 689
rect 52 665 171 669
rect 223 718 227 722
rect 223 703 227 707
rect 223 688 227 692
rect 223 673 227 677
rect 259 746 398 750
rect 402 746 411 770
rect 259 716 398 720
rect 402 696 411 720
rect 32 632 36 636
rect 1 521 5 625
rect 14 621 28 625
rect 14 584 18 618
rect 24 584 28 618
rect 39 619 173 623
rect 39 609 173 613
rect 39 599 173 603
rect 39 589 173 593
rect 279 665 398 669
rect 402 665 411 689
rect 414 641 418 645
rect 421 648 425 987
rect 414 634 418 638
rect 275 614 434 618
rect 275 604 434 608
rect 24 556 28 560
rect 24 546 28 550
rect 50 556 54 560
rect 50 546 54 550
rect 68 556 72 560
rect 68 546 72 550
rect 86 556 90 560
rect 86 546 90 550
rect 104 556 108 560
rect 104 546 108 550
rect 122 556 126 560
rect 122 546 126 550
rect 131 546 135 550
rect 2 480 6 484
rect 7 485 11 489
rect 28 503 32 512
rect 2 470 6 474
rect 149 546 153 550
rect 41 521 55 525
rect 35 495 44 499
rect 41 484 45 488
rect 51 484 55 488
rect 68 521 92 525
rect 105 521 129 525
rect 132 511 141 515
rect 95 503 104 507
rect 92 495 101 499
rect 64 484 68 488
rect 74 484 78 488
rect 84 484 88 488
rect 105 484 109 488
rect 115 484 119 488
rect 125 484 129 488
rect 138 503 147 507
rect 150 495 159 499
rect 167 494 171 503
rect 150 484 154 488
rect 160 484 164 488
rect 24 467 28 471
rect 2 460 6 464
rect 2 450 6 454
rect 2 440 6 444
rect 2 430 6 434
rect 2 420 6 424
rect 24 457 28 461
rect 24 447 28 451
rect 24 437 28 441
rect 24 427 28 431
rect 50 467 54 471
rect 50 457 54 461
rect 50 447 54 451
rect 50 437 54 441
rect 50 427 54 431
rect 68 467 72 471
rect 68 457 72 461
rect 68 447 72 451
rect 68 437 72 441
rect 68 427 72 431
rect 86 467 90 471
rect 86 457 90 461
rect 86 447 90 451
rect 86 437 90 441
rect 86 427 90 431
rect 104 467 108 471
rect 104 457 108 461
rect 104 447 108 451
rect 104 437 108 441
rect 104 427 108 431
rect 122 467 126 471
rect 122 457 126 461
rect 122 447 126 451
rect 122 437 126 441
rect 122 427 126 431
rect 149 462 153 466
rect 184 556 188 560
rect 184 546 188 550
rect 211 556 215 560
rect 211 546 215 550
rect 188 526 192 530
rect 190 511 199 515
rect 167 462 171 466
rect 185 467 189 471
rect 215 526 219 530
rect 222 494 226 503
rect 185 457 189 461
rect 185 447 189 451
rect 185 437 189 441
rect 185 427 189 431
rect 2 410 6 414
rect 2 400 6 404
rect 2 390 6 394
rect 212 467 216 471
rect 212 457 216 461
rect 212 447 216 451
rect 212 437 216 441
rect 212 427 216 431
rect 20 407 29 411
rect 20 397 29 401
rect 20 387 29 391
rect 32 407 36 411
rect 25 31 29 360
rect 32 365 36 374
rect 20 21 39 25
rect 49 407 53 411
rect 49 398 223 402
rect 49 387 173 391
rect 278 576 317 580
rect 276 566 325 570
rect 276 556 325 560
rect 276 546 325 550
rect 339 556 343 560
rect 339 546 343 550
rect 276 536 325 540
rect 276 521 345 525
rect 357 556 361 560
rect 357 546 361 550
rect 375 556 379 560
rect 375 546 379 550
rect 393 556 397 560
rect 393 546 397 550
rect 356 521 365 525
rect 348 501 352 510
rect 276 478 325 482
rect 276 468 325 472
rect 276 458 325 462
rect 276 448 325 452
rect 276 438 325 442
rect 276 428 325 432
rect 49 320 53 344
rect 57 340 171 344
rect 276 418 325 422
rect 276 408 325 412
rect 339 467 343 471
rect 339 457 343 461
rect 339 447 343 451
rect 339 437 343 441
rect 339 427 343 431
rect 355 483 359 487
rect 375 521 399 525
rect 380 483 384 487
rect 390 483 394 487
rect 357 467 361 471
rect 357 457 361 461
rect 357 447 361 451
rect 357 437 361 441
rect 357 427 361 431
rect 375 467 379 471
rect 375 457 379 461
rect 375 447 379 451
rect 375 437 379 441
rect 375 422 379 431
rect 393 467 397 471
rect 393 457 397 461
rect 393 447 397 451
rect 393 437 397 441
rect 393 427 397 431
rect 411 556 415 560
rect 411 546 415 550
rect 429 556 433 560
rect 429 546 433 550
rect 409 521 418 525
rect 429 521 438 525
rect 445 521 449 625
rect 421 501 425 510
rect 409 483 413 487
rect 434 485 438 489
rect 411 462 415 466
rect 411 452 415 456
rect 411 442 415 446
rect 411 432 415 436
rect 276 398 360 402
rect 276 387 395 391
rect 49 288 53 312
rect 223 333 227 337
rect 223 318 227 322
rect 277 340 396 344
rect 57 288 181 292
rect 49 238 53 262
rect 57 258 181 262
rect 49 207 53 231
rect 57 207 181 211
rect 49 157 53 181
rect 57 177 181 181
rect 223 260 227 264
rect 223 245 227 249
rect 223 230 227 234
rect 223 215 227 219
rect 267 288 396 292
rect 267 258 396 262
rect 267 207 396 211
rect 267 177 396 181
rect 49 126 53 150
rect 57 126 181 130
rect 49 76 53 100
rect 57 96 181 100
rect 223 163 227 167
rect 223 148 227 152
rect 223 133 227 137
rect 223 118 227 122
rect 267 126 396 130
rect 267 96 396 100
rect 49 45 53 69
rect 57 45 171 49
rect 50 27 169 31
rect 50 17 169 21
rect 223 67 227 71
rect 223 52 227 56
rect 178 15 272 29
rect 277 45 396 49
rect 280 27 399 31
rect 280 17 399 21
rect 11 9 20 13
rect 38 9 47 13
rect 395 9 404 13
rect 434 408 438 477
rect 414 397 438 401
rect 414 387 438 391
rect 445 385 449 489
rect 414 365 418 374
rect 421 31 425 360
rect 431 31 435 360
rect 416 20 435 24
rect 408 9 417 13
<< metal2 >>
rect 30 1495 420 1500
rect 30 1114 34 1495
rect 415 1114 420 1495
rect 30 1110 420 1114
rect 0 987 450 1010
rect 0 648 25 987
rect 29 986 421 987
rect 29 982 40 986
rect 174 982 421 986
rect 29 981 421 982
rect 29 977 280 981
rect 409 977 421 981
rect 29 964 421 977
rect 29 940 39 964
rect 48 960 52 964
rect 171 960 284 964
rect 398 960 402 964
rect 48 940 402 960
rect 411 940 421 964
rect 29 932 421 940
rect 29 908 39 932
rect 48 920 402 932
rect 48 916 223 920
rect 227 916 402 920
rect 48 912 402 916
rect 48 908 52 912
rect 191 908 264 912
rect 398 908 402 912
rect 411 908 421 932
rect 29 905 421 908
rect 29 901 223 905
rect 227 901 421 905
rect 29 890 421 901
rect 29 886 223 890
rect 227 886 421 890
rect 29 882 421 886
rect 29 858 39 882
rect 48 878 52 882
rect 191 878 264 882
rect 398 878 402 882
rect 48 875 402 878
rect 48 871 223 875
rect 227 871 402 875
rect 48 858 402 871
rect 411 858 421 882
rect 29 851 421 858
rect 29 827 39 851
rect 48 831 402 851
rect 48 827 52 831
rect 191 829 259 831
rect 191 827 223 829
rect 29 825 223 827
rect 227 827 259 829
rect 398 827 402 831
rect 411 827 421 851
rect 227 825 421 827
rect 29 814 421 825
rect 29 810 223 814
rect 227 810 421 814
rect 29 801 421 810
rect 29 777 39 801
rect 48 797 52 801
rect 191 799 259 801
rect 191 797 223 799
rect 48 795 223 797
rect 227 797 259 799
rect 398 797 402 801
rect 227 795 402 797
rect 48 784 402 795
rect 48 780 223 784
rect 227 780 402 784
rect 48 777 402 780
rect 411 777 421 801
rect 29 770 421 777
rect 29 746 39 770
rect 48 750 402 770
rect 48 746 52 750
rect 191 746 259 750
rect 398 746 402 750
rect 411 746 421 770
rect 29 722 421 746
rect 29 720 223 722
rect 29 696 39 720
rect 48 716 52 720
rect 191 718 223 720
rect 227 720 421 722
rect 227 718 259 720
rect 191 716 259 718
rect 398 716 402 720
rect 48 707 402 716
rect 48 703 223 707
rect 227 703 402 707
rect 48 696 402 703
rect 411 696 421 720
rect 29 692 421 696
rect 29 689 223 692
rect 29 665 39 689
rect 48 688 223 689
rect 227 689 421 692
rect 227 688 402 689
rect 48 677 402 688
rect 48 673 223 677
rect 227 673 402 677
rect 48 669 402 673
rect 48 665 52 669
rect 171 665 279 669
rect 398 665 402 669
rect 411 665 421 689
rect 29 649 421 665
rect 39 648 411 649
rect 425 648 450 987
rect 36 641 414 644
rect 32 638 418 641
rect 32 636 414 638
rect 36 634 414 636
rect 36 632 418 634
rect 0 625 450 626
rect 0 521 1 625
rect 5 621 14 625
rect 28 623 445 625
rect 28 621 39 623
rect 5 619 39 621
rect 173 619 445 623
rect 5 618 445 619
rect 5 584 14 618
rect 18 584 24 618
rect 28 614 275 618
rect 434 614 445 618
rect 28 613 445 614
rect 28 609 39 613
rect 173 609 445 613
rect 28 608 445 609
rect 28 604 275 608
rect 434 604 445 608
rect 28 603 445 604
rect 28 599 39 603
rect 173 599 445 603
rect 28 593 445 599
rect 28 589 39 593
rect 173 589 445 593
rect 28 584 445 589
rect 5 580 445 584
rect 5 576 278 580
rect 317 576 445 580
rect 5 570 445 576
rect 5 566 276 570
rect 325 566 445 570
rect 5 560 445 566
rect 5 556 24 560
rect 28 556 50 560
rect 54 556 68 560
rect 72 556 86 560
rect 90 556 104 560
rect 108 556 122 560
rect 126 556 184 560
rect 188 556 211 560
rect 215 556 276 560
rect 325 556 339 560
rect 343 556 357 560
rect 361 556 375 560
rect 379 556 393 560
rect 397 556 411 560
rect 415 556 429 560
rect 433 556 445 560
rect 5 554 445 556
rect 5 550 127 554
rect 157 550 445 554
rect 5 546 24 550
rect 28 546 50 550
rect 54 546 68 550
rect 72 546 86 550
rect 90 546 104 550
rect 108 546 122 550
rect 126 546 127 550
rect 135 546 149 550
rect 157 546 184 550
rect 188 546 211 550
rect 215 546 276 550
rect 325 546 339 550
rect 343 546 357 550
rect 361 546 375 550
rect 379 546 393 550
rect 397 546 411 550
rect 415 546 429 550
rect 433 546 445 550
rect 5 542 127 546
rect 157 542 445 546
rect 5 540 445 542
rect 5 536 276 540
rect 325 536 445 540
rect 5 530 445 536
rect 5 526 188 530
rect 192 526 215 530
rect 219 526 445 530
rect 5 525 445 526
rect 5 521 41 525
rect 55 521 68 525
rect 92 521 105 525
rect 129 521 276 525
rect 345 521 356 525
rect 365 521 375 525
rect 399 521 409 525
rect 418 521 429 525
rect 438 521 445 525
rect 449 521 450 625
rect 141 511 190 515
rect 32 503 95 507
rect 104 503 138 507
rect 44 495 92 499
rect 101 495 150 499
rect 171 494 222 503
rect 352 501 421 510
rect 0 485 7 489
rect 11 488 434 489
rect 11 485 41 488
rect 0 484 41 485
rect 45 484 51 488
rect 55 484 64 488
rect 68 484 74 488
rect 78 484 84 488
rect 88 484 105 488
rect 109 484 115 488
rect 119 484 125 488
rect 129 484 150 488
rect 154 484 160 488
rect 164 487 434 488
rect 164 484 355 487
rect 0 480 2 484
rect 6 483 355 484
rect 359 483 380 487
rect 384 483 390 487
rect 394 483 409 487
rect 413 485 434 487
rect 438 485 445 489
rect 413 483 445 485
rect 6 482 445 483
rect 6 480 276 482
rect 0 478 276 480
rect 325 478 445 482
rect 0 477 445 478
rect 0 474 434 477
rect 0 470 2 474
rect 6 472 434 474
rect 6 471 276 472
rect 6 470 24 471
rect 0 467 24 470
rect 28 467 50 471
rect 54 467 68 471
rect 72 467 86 471
rect 90 467 104 471
rect 108 467 122 471
rect 126 470 185 471
rect 126 467 145 470
rect 0 464 145 467
rect 175 467 185 470
rect 189 467 212 471
rect 216 468 276 471
rect 325 471 434 472
rect 325 468 339 471
rect 216 467 339 468
rect 343 467 357 471
rect 361 467 375 471
rect 379 467 393 471
rect 397 467 434 471
rect 175 466 434 467
rect 0 460 2 464
rect 6 461 145 464
rect 153 462 167 466
rect 175 462 411 466
rect 415 462 434 466
rect 6 460 24 461
rect 0 457 24 460
rect 28 457 50 461
rect 54 457 68 461
rect 72 457 86 461
rect 90 457 104 461
rect 108 457 122 461
rect 126 458 145 461
rect 175 461 276 462
rect 175 458 185 461
rect 126 457 185 458
rect 189 457 212 461
rect 216 458 276 461
rect 325 461 434 462
rect 325 458 339 461
rect 216 457 339 458
rect 343 457 357 461
rect 361 457 375 461
rect 379 457 393 461
rect 397 457 434 461
rect 0 456 434 457
rect 0 454 411 456
rect 0 450 2 454
rect 6 452 411 454
rect 415 452 434 456
rect 6 451 276 452
rect 6 450 24 451
rect 0 447 24 450
rect 28 447 50 451
rect 54 447 68 451
rect 72 447 86 451
rect 90 447 104 451
rect 108 447 122 451
rect 126 447 185 451
rect 189 447 212 451
rect 216 448 276 451
rect 325 451 434 452
rect 325 448 339 451
rect 216 447 339 448
rect 343 447 357 451
rect 361 447 375 451
rect 379 447 393 451
rect 397 447 434 451
rect 0 446 434 447
rect 0 444 411 446
rect 0 440 2 444
rect 6 442 411 444
rect 415 442 434 446
rect 6 441 276 442
rect 6 440 24 441
rect 0 437 24 440
rect 28 437 50 441
rect 54 437 68 441
rect 72 437 86 441
rect 90 437 104 441
rect 108 437 122 441
rect 126 437 185 441
rect 189 437 212 441
rect 216 438 276 441
rect 325 441 434 442
rect 325 438 339 441
rect 216 437 339 438
rect 343 437 357 441
rect 361 437 375 441
rect 379 437 393 441
rect 397 437 434 441
rect 0 436 434 437
rect 0 434 411 436
rect 0 430 2 434
rect 6 432 411 434
rect 415 432 434 436
rect 6 431 276 432
rect 6 430 24 431
rect 0 427 24 430
rect 28 427 50 431
rect 54 427 68 431
rect 72 427 86 431
rect 90 427 104 431
rect 108 427 122 431
rect 126 427 185 431
rect 189 427 212 431
rect 216 428 276 431
rect 325 431 434 432
rect 325 428 339 431
rect 216 427 339 428
rect 343 427 357 431
rect 361 427 375 431
rect 0 424 375 427
rect 0 420 2 424
rect 6 422 375 424
rect 379 427 393 431
rect 397 427 434 431
rect 379 422 434 427
rect 6 420 276 422
rect 0 418 276 420
rect 325 418 434 422
rect 0 415 434 418
rect 0 414 28 415
rect 0 410 2 414
rect 6 411 28 414
rect 57 412 434 415
rect 6 410 20 411
rect 0 407 20 410
rect 36 407 49 411
rect 57 408 276 412
rect 325 408 434 412
rect 438 408 445 477
rect 0 404 29 407
rect 0 400 2 404
rect 6 403 29 404
rect 57 403 445 408
rect 6 402 445 403
rect 6 401 49 402
rect 6 400 20 401
rect 0 397 20 400
rect 29 398 49 401
rect 223 398 276 402
rect 360 401 445 402
rect 360 398 414 401
rect 29 397 414 398
rect 438 397 445 401
rect 0 394 445 397
rect 0 390 2 394
rect 6 391 445 394
rect 6 390 20 391
rect 0 387 20 390
rect 29 387 49 391
rect 173 387 276 391
rect 395 387 414 391
rect 438 387 445 391
rect 0 386 445 387
rect 0 384 49 386
rect 173 385 445 386
rect 449 385 450 489
rect 173 384 450 385
rect 413 383 440 384
rect 36 366 414 374
rect 0 361 29 362
rect 39 361 411 362
rect 421 361 450 362
rect 0 360 450 361
rect 0 31 25 360
rect 29 344 421 360
rect 29 320 49 344
rect 53 340 57 344
rect 171 340 277 344
rect 396 340 421 344
rect 53 337 421 340
rect 53 333 223 337
rect 227 333 421 337
rect 53 322 421 333
rect 53 320 223 322
rect 29 318 223 320
rect 227 318 421 322
rect 29 312 421 318
rect 29 288 49 312
rect 53 292 421 312
rect 53 288 57 292
rect 181 288 267 292
rect 396 288 421 292
rect 29 264 421 288
rect 29 262 223 264
rect 29 238 49 262
rect 53 258 57 262
rect 181 260 223 262
rect 227 262 421 264
rect 227 260 267 262
rect 181 258 267 260
rect 396 258 421 262
rect 53 249 421 258
rect 53 245 223 249
rect 227 245 421 249
rect 53 238 421 245
rect 29 234 421 238
rect 29 231 223 234
rect 29 207 49 231
rect 53 230 223 231
rect 227 230 421 234
rect 53 219 421 230
rect 53 215 223 219
rect 227 215 421 219
rect 53 211 421 215
rect 53 207 57 211
rect 181 207 267 211
rect 396 207 421 211
rect 29 181 421 207
rect 29 157 49 181
rect 53 177 57 181
rect 181 177 267 181
rect 396 177 421 181
rect 53 167 421 177
rect 53 163 223 167
rect 227 163 421 167
rect 53 157 421 163
rect 29 152 421 157
rect 29 150 223 152
rect 29 126 49 150
rect 53 148 223 150
rect 227 148 421 152
rect 53 137 421 148
rect 53 133 223 137
rect 227 133 421 137
rect 53 130 421 133
rect 53 126 57 130
rect 181 126 267 130
rect 396 126 421 130
rect 29 122 421 126
rect 29 118 223 122
rect 227 118 421 122
rect 29 100 421 118
rect 29 76 49 100
rect 53 96 57 100
rect 181 96 267 100
rect 396 96 421 100
rect 53 76 421 96
rect 29 71 421 76
rect 29 69 223 71
rect 29 45 49 69
rect 53 67 223 69
rect 227 67 421 71
rect 53 56 421 67
rect 53 52 223 56
rect 227 52 421 56
rect 53 49 421 52
rect 53 45 57 49
rect 171 45 277 49
rect 396 45 421 49
rect 29 34 421 45
rect 29 31 172 34
rect 0 27 50 31
rect 169 27 172 31
rect 278 31 421 34
rect 425 31 431 360
rect 435 31 450 360
rect 0 25 172 27
rect 0 21 20 25
rect 39 21 172 25
rect 0 17 50 21
rect 169 17 172 21
rect 0 0 7 17
rect 11 0 20 9
rect 24 0 34 17
rect 38 0 47 9
rect 51 0 172 17
rect 177 15 178 29
rect 272 15 273 29
rect 177 0 273 15
rect 278 27 280 31
rect 399 27 450 31
rect 278 24 450 27
rect 278 21 416 24
rect 278 17 280 21
rect 399 20 416 21
rect 435 20 450 24
rect 399 17 450 20
rect 278 0 391 17
rect 395 0 404 9
rect 408 0 417 9
rect 421 0 450 17
<< pad >>
rect 34 1114 415 1495
<< pseudo_rpoly >>
rect 236 599 429 600
rect 236 586 429 587
<< rpoly >>
rect 236 587 429 599
<< m2p >>
rect 13 -2 17 2
rect 41 -2 45 2
rect 411 -2 415 2
<< m4p >>
rect 211 1330 222 1342
<< labels >>
rlabel metal2 413 0 413 0 8 DI
rlabel metal2 43 0 43 0 8 DO
rlabel metal2 214 812 214 812 6 Vdd2
rlabel metal2 199 185 199 185 6 Gnd2
rlabel metal2 15 0 15 0 8 OEN
rlabel metal2 243 444 243 444 6 Vdd
rlabel metal2 243 581 243 581 6 Gnd
rlabel m4p 216 1336 216 1336 1 YPAD
<< end >>

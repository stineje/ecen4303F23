magic
tech scmos
timestamp 1069013294
<< nwell >>
rect -8 48 80 105
<< ntransistor >>
rect 7 6 9 26
rect 15 6 17 26
rect 23 6 25 26
rect 31 6 33 26
rect 39 6 41 26
rect 47 6 49 26
rect 55 6 57 26
rect 63 6 65 26
<< ptransistor >>
rect 7 54 9 94
rect 15 54 17 94
rect 23 54 25 94
rect 31 54 33 94
rect 39 54 41 94
rect 47 54 49 94
rect 55 54 57 94
rect 63 54 65 94
<< ndiffusion >>
rect 6 6 7 26
rect 9 6 10 26
rect 14 6 15 26
rect 17 6 18 26
rect 22 6 23 26
rect 25 6 26 26
rect 30 6 31 26
rect 33 6 34 26
rect 38 6 39 26
rect 41 6 42 26
rect 46 6 47 26
rect 49 6 50 26
rect 54 6 55 26
rect 57 6 58 26
rect 62 6 63 26
rect 65 6 66 26
<< pdiffusion >>
rect 6 54 7 94
rect 9 54 10 94
rect 14 54 15 94
rect 17 54 18 94
rect 22 54 23 94
rect 25 54 26 94
rect 30 54 31 94
rect 33 54 34 94
rect 38 54 39 94
rect 41 54 42 94
rect 46 54 47 94
rect 49 54 50 94
rect 54 54 55 94
rect 57 54 58 94
rect 62 54 63 94
rect 65 54 66 94
<< ndcontact >>
rect 2 6 6 26
rect 10 6 14 26
rect 18 6 22 26
rect 26 6 30 26
rect 34 6 38 26
rect 42 6 46 26
rect 50 6 54 26
rect 58 6 62 26
rect 66 6 70 26
<< pdcontact >>
rect 2 54 6 94
rect 10 54 14 94
rect 18 54 22 94
rect 26 54 30 94
rect 34 54 38 94
rect 42 54 46 94
rect 50 54 54 94
rect 58 54 62 94
rect 66 54 70 94
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
rect 46 -2 50 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
rect 46 98 50 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 31 94 33 96
rect 39 94 41 96
rect 47 94 49 96
rect 55 94 57 96
rect 63 94 65 96
rect 7 40 9 54
rect 15 40 17 54
rect 11 36 17 40
rect 7 26 9 36
rect 15 26 17 36
rect 23 40 25 54
rect 31 40 33 54
rect 23 36 24 40
rect 28 36 33 40
rect 23 26 25 36
rect 31 26 33 36
rect 39 26 41 54
rect 47 40 49 54
rect 55 40 57 54
rect 63 40 65 54
rect 45 36 49 40
rect 54 36 58 40
rect 62 36 65 40
rect 47 26 49 36
rect 55 26 57 36
rect 63 26 65 36
rect 7 4 9 6
rect 15 4 17 6
rect 23 4 25 6
rect 31 4 33 6
rect 39 4 41 6
rect 47 4 49 6
rect 55 4 57 6
rect 63 4 65 6
<< polycontact >>
rect 7 36 11 40
rect 24 36 28 40
rect 41 36 45 40
rect 58 36 62 40
<< metal1 >>
rect -2 102 74 103
rect 2 98 14 102
rect 18 98 30 102
rect 34 98 46 102
rect 50 98 74 102
rect -2 97 74 98
rect 2 94 6 97
rect 18 94 22 97
rect 34 94 38 97
rect 50 94 54 97
rect 66 94 70 97
rect 10 51 14 54
rect 26 51 30 54
rect 42 51 46 54
rect 58 51 62 54
rect 10 47 19 51
rect 26 47 37 51
rect 42 47 53 51
rect 58 47 70 51
rect 15 40 19 47
rect 33 40 37 47
rect 49 40 53 47
rect 2 36 7 40
rect 15 36 24 40
rect 33 36 41 40
rect 49 36 58 40
rect 2 33 6 36
rect 15 33 19 36
rect 33 33 37 36
rect 49 33 53 36
rect 66 33 70 47
rect 10 29 19 33
rect 26 29 37 33
rect 42 29 53 33
rect 58 29 70 33
rect 10 26 14 29
rect 26 26 30 29
rect 42 26 46 29
rect 58 26 62 29
rect 2 3 6 6
rect 18 3 22 6
rect 34 3 38 6
rect 50 3 54 6
rect 66 3 70 6
rect -2 2 74 3
rect 2 -2 14 2
rect 18 -2 30 2
rect 34 -2 46 2
rect 50 -2 74 2
rect -2 -3 74 -2
<< m1p >>
rect 66 43 70 47
rect 2 33 6 37
<< labels >>
<< end >>

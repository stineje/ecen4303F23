module sram (A, D, Q, w, e);
input  [7:0] A,D ;
output [7:0] Q ;
input  w,e ;
endmodule

magic
tech scmos
timestamp 1052875792
use PADFC padfc_0
timestamp 949001400
transform 1 0 -305 0 1 -2
box 327 -3 1003 673
use PADGND padgnd_0
timestamp 1048632339
transform 1 0 724 0 1 -3
box -3 -3 303 1000
use PADINC padinc_0
timestamp 1052875792
transform 1 0 1054 0 1 -3
box -6 -3 303 1000
use PADOUT padout_0
timestamp 1052875792
transform 1 0 1382 0 1 8
box -6 -3 303 1000
use PADNC padnc_0
timestamp 1022363748
transform 1 0 1710 0 1 11
box -3 -3 303 1000
use PADVDD padvdd_0
timestamp 1048632506
transform 1 0 2034 0 1 12
box -3 -4 303 999
use PADINOUT PADINOUT_0
timestamp 1052875792
transform 1 0 2367 0 1 9
box -6 -3 303 1000
<< end >>

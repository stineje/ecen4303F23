magic
tech scmos
timestamp 1084294400
<< nwell >>
rect 20 740 280 1000
rect 17 429 283 653
rect -3 249 303 330
rect -3 11 11 249
rect 289 11 303 249
rect -3 -3 303 11
<< pwell >>
rect -3 656 303 673
rect -3 426 14 656
rect 286 426 303 656
rect -3 340 303 426
rect 11 11 289 249
<< psubstratepdiff >>
rect 0 668 300 670
rect 0 664 2 668
rect 166 664 169 668
rect 298 664 300 668
rect 0 662 300 664
rect 0 423 2 662
rect 6 659 294 662
rect 6 423 11 659
rect 289 423 294 659
rect 298 423 300 662
rect 0 413 300 423
rect 0 409 3 413
rect 297 409 300 413
rect 0 403 300 409
rect 0 399 3 403
rect 297 399 300 403
rect 0 393 300 399
rect 0 389 3 393
rect 297 389 300 393
rect 0 383 300 389
rect 0 379 3 383
rect 297 379 300 383
rect 0 373 300 379
rect 0 369 3 373
rect 297 369 300 373
rect 0 363 300 369
rect 0 359 3 363
rect 297 359 300 363
rect 0 353 300 359
rect 0 349 3 353
rect 297 349 300 353
rect 0 343 300 349
rect 14 245 286 246
rect 14 231 16 245
rect 285 231 286 245
rect 14 224 286 231
rect 14 220 16 224
rect 285 220 286 224
rect 14 214 286 220
rect 14 210 16 214
rect 285 210 286 214
rect 14 204 286 210
rect 14 200 16 204
rect 285 200 286 204
rect 14 194 286 200
rect 14 190 16 194
rect 285 190 286 194
rect 14 184 286 190
rect 14 180 16 184
rect 285 180 286 184
rect 14 174 286 180
rect 14 170 16 174
rect 285 170 286 174
rect 14 164 286 170
rect 14 160 16 164
rect 285 160 286 164
rect 14 154 286 160
rect 14 150 16 154
rect 285 150 286 154
rect 14 144 286 150
rect 14 140 16 144
rect 285 140 286 144
rect 14 134 286 140
rect 14 130 16 134
rect 285 130 286 134
rect 14 124 286 130
rect 14 120 16 124
rect 285 120 286 124
rect 14 114 286 120
rect 14 110 16 114
rect 285 110 286 114
rect 14 104 286 110
rect 14 100 16 104
rect 285 100 286 104
rect 14 94 286 100
rect 14 90 16 94
rect 285 90 286 94
rect 14 84 286 90
rect 14 80 16 84
rect 285 80 286 84
rect 14 74 286 80
rect 14 70 16 74
rect 285 70 286 74
rect 14 64 286 70
rect 14 60 16 64
rect 285 60 286 64
rect 14 54 286 60
rect 14 50 16 54
rect 285 50 286 54
rect 14 44 286 50
rect 14 40 16 44
rect 285 40 286 44
rect 14 34 286 40
rect 14 30 16 34
rect 285 30 286 34
rect 14 24 286 30
rect 14 20 16 24
rect 285 20 286 24
rect 14 14 286 20
<< nsubstratendiff >>
rect 20 649 280 650
rect 20 645 23 649
rect 277 645 280 649
rect 20 639 280 645
rect 20 635 23 639
rect 277 635 280 639
rect 20 629 280 635
rect 20 625 23 629
rect 277 625 280 629
rect 20 619 280 625
rect 20 615 23 619
rect 277 615 280 619
rect 20 609 280 615
rect 20 605 23 609
rect 277 605 280 609
rect 20 599 280 605
rect 20 595 23 599
rect 277 595 280 599
rect 20 589 280 595
rect 20 585 23 589
rect 277 585 280 589
rect 20 579 280 585
rect 20 575 23 579
rect 277 575 280 579
rect 20 569 280 575
rect 20 565 23 569
rect 277 565 280 569
rect 20 559 280 565
rect 20 555 23 559
rect 277 555 280 559
rect 20 549 280 555
rect 20 545 23 549
rect 277 545 280 549
rect 20 539 280 545
rect 20 535 23 539
rect 277 535 280 539
rect 20 529 280 535
rect 20 525 23 529
rect 277 525 280 529
rect 20 519 280 525
rect 20 515 23 519
rect 277 515 280 519
rect 20 509 280 515
rect 20 505 23 509
rect 277 505 280 509
rect 20 499 280 505
rect 20 495 23 499
rect 277 495 280 499
rect 20 489 280 495
rect 20 485 23 489
rect 277 485 280 489
rect 20 479 280 485
rect 20 475 23 479
rect 277 475 280 479
rect 20 469 280 475
rect 20 465 23 469
rect 277 465 280 469
rect 20 459 280 465
rect 20 455 23 459
rect 277 455 280 459
rect 20 449 280 455
rect 20 445 23 449
rect 277 445 280 449
rect 20 438 280 445
rect 20 434 23 438
rect 277 434 280 438
rect 20 432 280 434
rect 0 323 300 327
rect 0 319 3 323
rect 297 319 300 323
rect 0 313 300 319
rect 0 309 3 313
rect 297 309 300 313
rect 0 303 300 309
rect 0 299 3 303
rect 297 299 300 303
rect 0 293 300 299
rect 0 289 3 293
rect 297 289 300 293
rect 0 283 300 289
rect 0 279 3 283
rect 297 279 300 283
rect 0 273 300 279
rect 0 269 3 273
rect 297 269 300 273
rect 0 263 300 269
rect 0 259 3 263
rect 297 259 300 263
rect 0 252 300 259
rect 0 251 8 252
rect 0 2 2 251
rect 6 8 8 251
rect 292 251 300 252
rect 292 8 294 251
rect 6 6 294 8
rect 6 2 8 6
rect 292 2 294 6
rect 298 2 300 251
rect 0 0 300 2
<< psubstratepcontact >>
rect 2 664 166 668
rect 169 664 298 668
rect 2 423 6 662
rect 294 423 298 662
rect 3 409 297 413
rect 3 399 297 403
rect 3 389 297 393
rect 3 379 297 383
rect 3 369 297 373
rect 3 359 297 363
rect 3 349 297 353
rect 16 231 285 245
rect 16 220 285 224
rect 16 210 285 214
rect 16 200 285 204
rect 16 190 285 194
rect 16 180 285 184
rect 16 170 285 174
rect 16 160 285 164
rect 16 150 285 154
rect 16 140 285 144
rect 16 130 285 134
rect 16 120 285 124
rect 16 110 285 114
rect 16 100 285 104
rect 16 90 285 94
rect 16 80 285 84
rect 16 70 285 74
rect 16 60 285 64
rect 16 50 285 54
rect 16 40 285 44
rect 16 30 285 34
rect 16 20 285 24
<< nsubstratencontact >>
rect 23 645 277 649
rect 23 635 277 639
rect 23 625 277 629
rect 23 615 277 619
rect 23 605 277 609
rect 23 595 277 599
rect 23 585 277 589
rect 23 575 277 579
rect 23 565 277 569
rect 23 555 277 559
rect 23 545 277 549
rect 23 535 277 539
rect 23 525 277 529
rect 23 515 277 519
rect 23 505 277 509
rect 23 495 277 499
rect 23 485 277 489
rect 23 475 277 479
rect 23 465 277 469
rect 23 455 277 459
rect 23 445 277 449
rect 23 434 277 438
rect 3 319 297 323
rect 3 309 297 313
rect 3 299 297 303
rect 3 289 297 293
rect 3 279 297 283
rect 3 269 297 273
rect 3 259 297 263
rect 2 2 6 251
rect 8 2 292 6
rect 294 2 298 251
<< metal1 >>
rect 20 997 280 1000
rect 20 743 23 997
rect 277 743 280 997
rect 20 740 280 743
rect 0 668 300 670
rect 0 664 2 668
rect 166 664 169 668
rect 298 664 300 668
rect 0 663 300 664
rect 0 662 7 663
rect 0 423 2 662
rect 6 423 7 662
rect 293 662 300 663
rect 21 645 23 649
rect 277 645 280 649
rect 21 644 280 645
rect 21 640 23 644
rect 277 640 280 644
rect 21 639 280 640
rect 21 635 23 639
rect 277 635 280 639
rect 21 634 280 635
rect 21 630 23 634
rect 277 630 280 634
rect 21 629 280 630
rect 21 625 23 629
rect 277 625 280 629
rect 21 624 280 625
rect 21 620 23 624
rect 277 620 280 624
rect 21 619 280 620
rect 21 615 23 619
rect 277 615 280 619
rect 21 614 280 615
rect 21 610 23 614
rect 277 610 280 614
rect 21 609 280 610
rect 21 605 23 609
rect 277 605 280 609
rect 21 604 280 605
rect 21 600 23 604
rect 277 600 280 604
rect 21 599 280 600
rect 21 595 23 599
rect 277 595 280 599
rect 21 594 280 595
rect 21 590 23 594
rect 277 590 280 594
rect 21 589 280 590
rect 21 585 23 589
rect 277 585 280 589
rect 21 584 280 585
rect 21 580 23 584
rect 277 580 280 584
rect 21 579 280 580
rect 21 575 23 579
rect 277 575 280 579
rect 21 574 280 575
rect 21 570 23 574
rect 277 570 280 574
rect 21 569 280 570
rect 21 565 23 569
rect 277 565 280 569
rect 21 564 280 565
rect 21 560 23 564
rect 277 560 280 564
rect 21 559 280 560
rect 21 555 23 559
rect 277 555 280 559
rect 21 554 280 555
rect 21 550 23 554
rect 277 550 280 554
rect 21 549 280 550
rect 21 545 23 549
rect 277 545 280 549
rect 21 544 280 545
rect 21 540 23 544
rect 277 540 280 544
rect 21 539 280 540
rect 21 535 23 539
rect 277 535 280 539
rect 21 534 280 535
rect 21 530 23 534
rect 277 530 280 534
rect 21 529 280 530
rect 21 525 23 529
rect 277 525 280 529
rect 21 524 280 525
rect 21 520 23 524
rect 277 520 280 524
rect 21 519 280 520
rect 21 515 23 519
rect 277 515 280 519
rect 21 514 280 515
rect 21 510 23 514
rect 277 510 280 514
rect 21 509 280 510
rect 21 505 23 509
rect 277 505 280 509
rect 21 504 280 505
rect 21 500 23 504
rect 277 500 280 504
rect 21 499 280 500
rect 21 495 23 499
rect 277 495 280 499
rect 21 494 280 495
rect 21 490 23 494
rect 277 490 280 494
rect 21 489 280 490
rect 21 485 23 489
rect 277 485 280 489
rect 21 484 280 485
rect 21 480 23 484
rect 277 480 280 484
rect 21 479 280 480
rect 21 475 23 479
rect 277 475 280 479
rect 21 474 280 475
rect 21 470 23 474
rect 277 470 280 474
rect 21 469 280 470
rect 21 465 23 469
rect 277 465 280 469
rect 21 464 280 465
rect 21 460 23 464
rect 277 460 280 464
rect 21 459 280 460
rect 21 455 23 459
rect 277 455 280 459
rect 21 454 280 455
rect 21 450 23 454
rect 277 450 280 454
rect 21 449 280 450
rect 21 445 23 449
rect 277 445 280 449
rect 21 444 280 445
rect 21 440 23 444
rect 277 440 280 444
rect 21 438 280 440
rect 21 434 23 438
rect 277 434 280 438
rect 21 433 280 434
rect 0 419 7 423
rect 293 423 294 662
rect 298 423 300 662
rect 293 419 300 423
rect 0 418 300 419
rect 0 414 3 418
rect 297 414 300 418
rect 0 413 300 414
rect 0 409 3 413
rect 297 409 300 413
rect 0 408 300 409
rect 0 404 3 408
rect 297 404 300 408
rect 0 403 300 404
rect 0 399 3 403
rect 297 399 300 403
rect 0 398 300 399
rect 0 394 3 398
rect 297 394 300 398
rect 0 393 300 394
rect 0 389 3 393
rect 297 389 300 393
rect 0 388 300 389
rect 0 384 3 388
rect 297 384 300 388
rect 0 383 300 384
rect 0 379 3 383
rect 297 379 300 383
rect 0 378 300 379
rect 0 374 3 378
rect 297 374 300 378
rect 0 373 300 374
rect 0 369 3 373
rect 297 369 300 373
rect 0 368 300 369
rect 0 364 3 368
rect 297 364 300 368
rect 0 363 300 364
rect 0 359 3 363
rect 297 359 300 363
rect 0 358 300 359
rect 0 354 3 358
rect 297 354 300 358
rect 0 353 300 354
rect 0 349 3 353
rect 297 349 300 353
rect 0 348 300 349
rect 0 344 3 348
rect 297 344 300 348
rect 0 323 300 326
rect 0 319 3 323
rect 297 319 300 323
rect 0 318 300 319
rect 0 314 3 318
rect 297 314 300 318
rect 0 313 300 314
rect 0 309 3 313
rect 297 309 300 313
rect 0 308 300 309
rect 0 304 3 308
rect 297 304 300 308
rect 0 303 300 304
rect 0 299 3 303
rect 297 299 300 303
rect 0 298 300 299
rect 0 294 3 298
rect 297 294 300 298
rect 0 293 300 294
rect 0 289 3 293
rect 297 289 300 293
rect 0 288 300 289
rect 0 284 3 288
rect 297 284 300 288
rect 0 283 300 284
rect 0 279 3 283
rect 297 279 300 283
rect 0 278 300 279
rect 0 274 3 278
rect 297 274 300 278
rect 0 273 300 274
rect 0 269 3 273
rect 297 269 300 273
rect 0 268 300 269
rect 0 264 3 268
rect 297 264 300 268
rect 0 263 300 264
rect 0 259 3 263
rect 297 259 300 263
rect 0 258 300 259
rect 0 254 3 258
rect 297 254 300 258
rect 0 253 300 254
rect 0 251 7 253
rect 0 2 2 251
rect 6 7 7 251
rect 293 251 300 253
rect 15 231 16 245
rect 15 229 285 231
rect 15 225 16 229
rect 285 225 286 229
rect 15 224 286 225
rect 15 220 16 224
rect 285 220 286 224
rect 15 219 286 220
rect 15 215 16 219
rect 285 215 286 219
rect 15 214 286 215
rect 15 210 16 214
rect 285 210 286 214
rect 15 209 286 210
rect 15 205 16 209
rect 285 205 286 209
rect 15 204 286 205
rect 15 200 16 204
rect 285 200 286 204
rect 15 199 286 200
rect 15 195 16 199
rect 285 195 286 199
rect 15 194 286 195
rect 15 190 16 194
rect 285 190 286 194
rect 15 189 286 190
rect 15 185 16 189
rect 285 185 286 189
rect 15 184 286 185
rect 15 180 16 184
rect 285 180 286 184
rect 15 179 286 180
rect 15 175 16 179
rect 285 175 286 179
rect 15 174 286 175
rect 15 170 16 174
rect 285 170 286 174
rect 15 169 286 170
rect 15 165 16 169
rect 285 165 286 169
rect 15 164 286 165
rect 15 160 16 164
rect 285 160 286 164
rect 15 159 286 160
rect 15 155 16 159
rect 285 155 286 159
rect 15 154 286 155
rect 15 150 16 154
rect 285 150 286 154
rect 15 149 286 150
rect 15 145 16 149
rect 285 145 286 149
rect 15 144 286 145
rect 15 140 16 144
rect 285 140 286 144
rect 15 139 286 140
rect 15 135 16 139
rect 285 135 286 139
rect 15 134 286 135
rect 15 130 16 134
rect 285 130 286 134
rect 15 129 286 130
rect 15 125 16 129
rect 285 125 286 129
rect 15 124 286 125
rect 15 120 16 124
rect 285 120 286 124
rect 15 119 286 120
rect 15 115 16 119
rect 285 115 286 119
rect 15 114 286 115
rect 15 110 16 114
rect 285 110 286 114
rect 15 109 286 110
rect 15 105 16 109
rect 285 105 286 109
rect 15 104 286 105
rect 15 100 16 104
rect 285 100 286 104
rect 15 99 286 100
rect 15 95 16 99
rect 285 95 286 99
rect 15 94 286 95
rect 15 90 16 94
rect 285 90 286 94
rect 15 89 286 90
rect 15 85 16 89
rect 285 85 286 89
rect 15 84 286 85
rect 15 80 16 84
rect 285 80 286 84
rect 15 79 286 80
rect 15 75 16 79
rect 285 75 286 79
rect 15 74 286 75
rect 15 70 16 74
rect 285 70 286 74
rect 15 69 286 70
rect 15 65 16 69
rect 285 65 286 69
rect 15 64 286 65
rect 15 60 16 64
rect 285 60 286 64
rect 15 59 286 60
rect 15 55 16 59
rect 285 55 286 59
rect 15 54 286 55
rect 15 50 16 54
rect 285 50 286 54
rect 15 49 286 50
rect 15 45 16 49
rect 285 45 286 49
rect 15 44 286 45
rect 15 40 16 44
rect 285 40 286 44
rect 15 39 286 40
rect 15 35 16 39
rect 285 35 286 39
rect 15 34 286 35
rect 15 30 16 34
rect 285 30 286 34
rect 15 29 286 30
rect 15 25 16 29
rect 285 25 286 29
rect 15 24 286 25
rect 15 20 16 24
rect 285 20 286 24
rect 15 19 286 20
rect 15 15 16 19
rect 285 15 286 19
rect 293 7 294 251
rect 6 6 294 7
rect 6 2 8 6
rect 292 2 294 6
rect 298 2 300 251
rect 0 1 300 2
<< m2contact >>
rect 23 640 277 644
rect 23 630 277 634
rect 23 620 277 624
rect 23 610 277 614
rect 23 600 277 604
rect 23 590 277 594
rect 23 580 277 584
rect 23 570 277 574
rect 23 560 277 564
rect 23 550 277 554
rect 23 540 277 544
rect 23 530 277 534
rect 23 520 277 524
rect 23 510 277 514
rect 23 500 277 504
rect 23 490 277 494
rect 23 480 277 484
rect 23 470 277 474
rect 23 460 277 464
rect 23 450 277 454
rect 23 440 277 444
rect 3 414 297 418
rect 3 404 297 408
rect 3 394 297 398
rect 3 384 297 388
rect 3 374 297 378
rect 3 364 297 368
rect 3 354 297 358
rect 3 344 297 348
rect 3 314 297 318
rect 3 304 297 308
rect 3 294 297 298
rect 3 284 297 288
rect 3 274 297 278
rect 3 264 297 268
rect 3 254 297 258
rect 16 225 285 229
rect 16 215 285 219
rect 16 205 285 209
rect 16 195 285 199
rect 16 185 285 189
rect 16 175 285 179
rect 16 165 285 169
rect 16 155 285 159
rect 16 145 285 149
rect 16 135 285 139
rect 16 125 285 129
rect 16 115 285 119
rect 16 105 285 109
rect 16 95 285 99
rect 16 85 285 89
rect 16 75 285 79
rect 16 65 285 69
rect 16 55 285 59
rect 16 45 285 49
rect 16 35 285 39
rect 16 25 285 29
rect 16 15 285 19
<< metal2 >>
rect 20 997 280 1000
rect 20 743 23 997
rect 277 743 280 997
rect 20 740 280 743
rect 0 644 300 670
rect 0 640 23 644
rect 277 640 300 644
rect 0 634 300 640
rect 0 630 23 634
rect 277 630 300 634
rect 0 624 300 630
rect 0 620 23 624
rect 277 620 300 624
rect 0 614 300 620
rect 0 610 23 614
rect 277 610 300 614
rect 0 604 300 610
rect 0 600 23 604
rect 277 600 300 604
rect 0 594 300 600
rect 0 590 23 594
rect 277 590 300 594
rect 0 584 300 590
rect 0 580 23 584
rect 277 580 300 584
rect 0 574 300 580
rect 0 570 23 574
rect 277 570 300 574
rect 0 564 300 570
rect 0 560 23 564
rect 277 560 300 564
rect 0 554 300 560
rect 0 550 23 554
rect 277 550 300 554
rect 0 544 300 550
rect 0 540 23 544
rect 277 540 300 544
rect 0 534 300 540
rect 0 530 23 534
rect 277 530 300 534
rect 0 524 300 530
rect 0 520 23 524
rect 277 520 300 524
rect 0 514 300 520
rect 0 510 23 514
rect 277 510 300 514
rect 0 504 300 510
rect 0 500 23 504
rect 277 500 300 504
rect 0 494 300 500
rect 0 490 23 494
rect 277 490 300 494
rect 0 484 300 490
rect 0 480 23 484
rect 277 480 300 484
rect 0 474 300 480
rect 0 470 23 474
rect 277 470 300 474
rect 0 464 300 470
rect 0 460 23 464
rect 277 460 300 464
rect 0 454 300 460
rect 0 450 23 454
rect 277 450 300 454
rect 0 444 300 450
rect 0 440 23 444
rect 277 440 300 444
rect 0 418 300 424
rect 0 414 3 418
rect 297 414 300 418
rect 0 408 300 414
rect 0 404 3 408
rect 297 404 300 408
rect 0 398 300 404
rect 0 394 3 398
rect 297 394 300 398
rect 0 388 300 394
rect 0 384 3 388
rect 297 384 300 388
rect 0 378 300 384
rect 0 374 3 378
rect 297 374 300 378
rect 0 368 300 374
rect 0 364 3 368
rect 297 364 300 368
rect 0 358 300 364
rect 0 354 3 358
rect 297 354 300 358
rect 0 348 300 354
rect 0 344 3 348
rect 297 344 300 348
rect 0 318 300 326
rect 0 314 3 318
rect 297 314 300 318
rect 0 308 300 314
rect 0 304 3 308
rect 297 304 300 308
rect 0 298 300 304
rect 0 294 3 298
rect 297 294 300 298
rect 0 288 300 294
rect 0 284 3 288
rect 297 284 300 288
rect 0 278 300 284
rect 0 274 3 278
rect 297 274 300 278
rect 0 268 300 274
rect 0 264 3 268
rect 297 264 300 268
rect 0 258 300 264
rect 0 254 3 258
rect 297 254 300 258
rect 0 246 300 254
rect 0 229 300 230
rect 0 225 16 229
rect 285 225 300 229
rect 0 219 300 225
rect 0 215 16 219
rect 285 215 300 219
rect 0 209 300 215
rect 0 205 16 209
rect 285 205 300 209
rect 0 199 300 205
rect 0 195 16 199
rect 285 195 300 199
rect 0 189 300 195
rect 0 185 16 189
rect 285 185 300 189
rect 0 179 300 185
rect 0 175 16 179
rect 285 175 300 179
rect 0 169 300 175
rect 0 165 16 169
rect 285 165 300 169
rect 0 159 300 165
rect 0 155 16 159
rect 285 155 300 159
rect 0 149 300 155
rect 0 145 16 149
rect 285 145 300 149
rect 0 139 300 145
rect 0 135 16 139
rect 285 135 300 139
rect 0 129 300 135
rect 0 125 16 129
rect 285 125 300 129
rect 0 119 300 125
rect 0 115 16 119
rect 285 115 300 119
rect 0 109 300 115
rect 0 105 16 109
rect 285 105 300 109
rect 0 99 300 105
rect 0 95 16 99
rect 285 95 300 99
rect 0 89 300 95
rect 0 85 16 89
rect 285 85 300 89
rect 0 79 300 85
rect 0 75 16 79
rect 285 75 300 79
rect 0 69 300 75
rect 0 65 16 69
rect 285 65 300 69
rect 0 59 300 65
rect 0 55 16 59
rect 285 55 300 59
rect 0 49 300 55
rect 0 45 16 49
rect 285 45 300 49
rect 0 39 300 45
rect 0 35 16 39
rect 285 35 300 39
rect 0 29 300 35
rect 0 25 16 29
rect 285 25 300 29
rect 0 19 300 25
rect 0 15 16 19
rect 285 15 300 19
rect 0 0 300 15
<< pad >>
rect 23 743 277 997
<< end >>

VERSION 5.3 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.05 ;

LAYER nwell
  TYPE	MASTERSLICE ;
END nwell

LAYER nactive
  TYPE	MASTERSLICE ;
END nactive

LAYER pactive
  TYPE	MASTERSLICE ;
END pactive

LAYER poly
  TYPE	MASTERSLICE ;
END poly

LAYER cc
  TYPE	CUT ;
  SPACING	0.45 ;
END cc

LAYER metal1
  TYPE		  ROUTING ;
  DIRECTION	  HORIZONTAL ;
  PITCH		  1.0  ;
  WIDTH		  0.3 ;
  SPACING	  0.3 ;
  RESISTANCE	  RPERSQ 0.08 ;
  CAPACITANCE	  CPERSQDIST 3.8e-05 ;
  EDGECAPACITANCE 8.0e-05 ;
  CURRENTDEN 0 ;
END metal1

LAYER via
  TYPE	CUT ;
  SPACING	0.3 ;
END via

LAYER metal2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.8  ;
  WIDTH		0.3 ;
  SPACING	0.3 ;
  RESISTANCE	RPERSQ 0.08 ;
  CAPACITANCE	CPERSQDIST 1.9e-05 ;
  EDGECAPACITANCE 6.0e-05 ;
  CURRENTDEN 0 ;
END metal2

LAYER via2
  TYPE	CUT ;
  SPACING	0.3 ;
END via2

LAYER metal3
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		1  ;
  WIDTH		0.3 ;
  SPACING	0.3 ;
  RESISTANCE	RPERSQ 0.08 ;
  CAPACITANCE	CPERSQDIST 1.3e-05 ;
  EDGECAPACITANCE 5.4e-05 ;
  CURRENTDEN 0 ;
END metal3

LAYER via3
  TYPE	CUT ;
  SPACING	0.4 ;
END via3

LAYER metal4
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.8  ;
  WIDTH		0.3 ;
  SPACING	0.3 ;
  RESISTANCE	RPERSQ 0.07 ;
  CAPACITANCE	CPERSQDIST 0.8e-05 ;
  EDGECAPACITANCE 4.1e-05 ;
  CURRENTDEN 0 ;
END metal4

LAYER via4
  TYPE	CUT ;
  SPACING	0.3 ;
END via4

LAYER metal5
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		1  ;
  WIDTH		0.3 ;
  SPACING	0.3 ;
  RESISTANCE	RPERSQ 0.07 ;
  CAPACITANCE	CPERSQDIST 0.8e-05 ;
  EDGECAPACITANCE 2.4e-05 ;
  CURRENTDEN 0 ;
END metal5

LAYER via5
  TYPE	CUT ;
  SPACING	0.4 ;
END via5

LAYER metal6
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		1.6 ;
  WIDTH		0.5 ;
  SPACING	0.5 ;
  RESISTANCE	RPERSQ 0.03 ;
  CAPACITANCE	CPERSQDIST 0.3e-05 ;
  EDGECAPACITANCE 2.0e-05 ;
  CURRENTDEN 0 ;
END metal6

VIA M6_M5 DEFAULT
  LAYER metal5 ;
    RECT -0.250 -0.250 0.250 0.250 ;
  LAYER via5 ;
    RECT -0.150 -0.150 0.150 0.150 ;
  LAYER metal6 ;
    RECT -0.250 -0.250 0.250 0.250 ;
END M6_M5

VIA M5_M4 DEFAULT
  LAYER metal4 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER via4 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER metal5 ;
    RECT -0.200 -0.200 0.200 0.200 ;
END M5_M4

VIA M4_M3 DEFAULT
  LAYER metal3 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER via3 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER metal4 ;
    RECT -0.200 -0.200 0.200 0.200 ;
END M4_M3

VIA M3_M2 DEFAULT
  LAYER metal2 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER via2 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER metal3 ;
    RECT -0.200 -0.200 0.200 0.200 ;
END M3_M2

VIA M2_M1 DEFAULT
  LAYER metal1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER via ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER metal2 ;
    RECT -0.200 -0.200 0.200 0.200 ;
END M2_M1


VIARULE viagen21 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.3 TO 60 ;
    OVERHANG 0.10 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 0.3 TO 60 ;
    OVERHANG 0.10 ;
    METALOVERHANG 0 ;
  LAYER via ;
    RECT -0.10 -0.10 0.10 0.10 ;
    SPACING 0.5 BY 0.5 ;
END viagen21

VIARULE viagen32 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.3 TO 60 ;
    OVERHANG 0.10 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 0.3 TO 60 ;
    OVERHANG 0.10 ;
    METALOVERHANG 0 ;
  LAYER via2 ;
    RECT -0.10 -0.10 0.10 0.10 ;
    SPACING 0.5 BY 0.5 ;
END viagen32

VIARULE viagen43 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.3 TO 60 ;
    OVERHANG 0.10 ;
    METALOVERHANG 0 ;
  LAYER metal4 ;
    DIRECTION VERTICAL ;
    WIDTH 0.3 TO 60 ;
    OVERHANG 0.10 ;
    METALOVERHANG 0 ;
  LAYER via3 ;
    RECT -0.10 -0.10 0.10 0.10 ;
    SPACING 0.6 BY 0.6 ;
END viagen43

VIARULE viagen54 GENERATE
  LAYER metal5 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.3 TO 60 ;
    OVERHANG 0.10 ;
    METALOVERHANG 0 ;
  LAYER metal4 ;
    DIRECTION VERTICAL ;
    WIDTH 0.3 TO 60 ;
    OVERHANG 0.10 ;
    METALOVERHANG 0 ;
  LAYER via4 ;
    RECT -0.10 -0.10 0.10 0.10 ;
    SPACING 0.5 BY 0.5 ;
END viagen54

VIARULE viagen65 GENERATE
  LAYER metal6 ;
    DIRECTION VERTICAL ;
    WIDTH 0.5 TO 60 ;
    OVERHANG 0.10 ;
    METALOVERHANG 0 ;
  LAYER metal5 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.5 TO 60 ;
    OVERHANG 0.10 ;
    METALOVERHANG 0 ;
  LAYER via5 ;
    RECT -0.15 -0.15 0.15 0.15 ;
    SPACING 0.7 BY 0.7 ;
END viagen65


VIARULE TURN1 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
  LAYER metal1 ;
    DIRECTION VERTICAL ;
END TURN1

VIARULE TURN2 GENERATE
  LAYER metal2 ;
    DIRECTION HORIZONTAL ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
END TURN2

VIARULE TURN3 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
  LAYER metal3 ;
    DIRECTION VERTICAL ;
END TURN3

VIARULE TURN4 GENERATE
  LAYER metal4 ;
    DIRECTION HORIZONTAL ;
  LAYER metal4 ;
    DIRECTION VERTICAL ;
END TURN4

VIARULE TURN5 GENERATE
  LAYER metal5 ;
    DIRECTION HORIZONTAL ;
  LAYER metal5 ;
    DIRECTION VERTICAL ;
END TURN5

VIARULE TURN6 GENERATE
  LAYER metal6 ;
    DIRECTION HORIZONTAL ;
  LAYER metal6 ;
    DIRECTION VERTICAL ;
END TURN6

SITE  core
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	0.800 BY 10.000 ;
END  core

END LIBRARY

magic
tech sky130A
timestamp 1605718197
<< psubdiff >>
rect -12 0 0 17
rect 17 0 29 17
<< psubdiffcont >>
rect 0 0 17 17
<< locali >>
rect -8 0 0 17
rect 17 0 25 17
<< end >>

magic
tech scmos
timestamp 1091055079
<< nwell >>
rect 30 1110 420 1500
<< hvnwell >>
rect 17 637 433 993
rect -3 376 453 493
rect -3 14 17 376
rect 433 14 453 376
rect -3 -3 453 14
<< hvpwell >>
rect -3 996 453 1013
rect -3 634 14 996
rect 436 634 453 996
rect -3 517 453 634
rect 17 14 433 376
<< hvptransistor >>
rect 38 965 213 968
rect 237 965 412 968
rect 38 904 213 907
rect 237 904 412 907
rect 38 883 213 886
rect 237 883 412 886
rect 38 823 213 826
rect 237 823 412 826
rect 38 802 213 805
rect 237 802 412 805
rect 38 742 213 745
rect 237 742 412 745
rect 38 721 213 724
rect 237 721 412 724
rect 38 661 213 664
rect 237 661 412 664
<< hvpdiffusion >>
rect 38 976 213 977
rect 38 972 41 976
rect 170 972 213 976
rect 38 968 213 972
rect 38 941 213 965
rect 38 937 61 941
rect 195 937 213 941
rect 38 935 213 937
rect 38 931 61 935
rect 195 931 213 935
rect 38 907 213 931
rect 237 976 412 977
rect 237 972 280 976
rect 409 972 412 976
rect 237 968 412 972
rect 237 941 412 965
rect 237 937 255 941
rect 389 937 412 941
rect 237 935 412 937
rect 237 931 255 935
rect 389 931 412 935
rect 237 907 412 931
rect 38 900 213 904
rect 38 896 46 900
rect 190 896 213 900
rect 38 894 213 896
rect 38 890 46 894
rect 190 890 213 894
rect 38 886 213 890
rect 237 900 412 904
rect 237 896 260 900
rect 404 896 412 900
rect 237 894 412 896
rect 237 890 260 894
rect 404 890 412 894
rect 237 886 412 890
rect 38 859 213 883
rect 38 850 61 859
rect 195 850 213 859
rect 38 826 213 850
rect 237 859 412 883
rect 237 850 255 859
rect 389 850 412 859
rect 237 826 412 850
rect 38 819 213 823
rect 38 815 46 819
rect 190 815 213 819
rect 38 813 213 815
rect 38 809 46 813
rect 190 809 213 813
rect 38 805 213 809
rect 38 778 213 802
rect 38 769 61 778
rect 195 769 213 778
rect 38 745 213 769
rect 237 819 412 823
rect 237 815 260 819
rect 404 815 412 819
rect 237 813 412 815
rect 237 809 260 813
rect 404 809 412 813
rect 237 805 412 809
rect 38 738 213 742
rect 38 734 46 738
rect 190 734 213 738
rect 38 732 213 734
rect 38 728 46 732
rect 190 728 213 732
rect 38 724 213 728
rect 237 778 412 802
rect 237 769 255 778
rect 389 769 412 778
rect 237 745 412 769
rect 237 738 412 742
rect 237 734 260 738
rect 404 734 412 738
rect 237 732 412 734
rect 237 728 260 732
rect 404 728 412 732
rect 237 724 412 728
rect 38 697 213 721
rect 38 688 61 697
rect 195 688 213 697
rect 38 664 213 688
rect 38 657 213 661
rect 38 653 41 657
rect 170 653 213 657
rect 38 652 213 653
rect 237 697 412 721
rect 237 688 255 697
rect 389 688 412 697
rect 237 664 412 688
rect 237 657 412 661
rect 237 653 280 657
rect 409 653 412 657
rect 237 652 412 653
<< hvpdcontact >>
rect 41 972 170 976
rect 61 937 195 941
rect 61 931 195 935
rect 280 972 409 976
rect 255 937 389 941
rect 255 931 389 935
rect 46 896 190 900
rect 46 890 190 894
rect 260 896 404 900
rect 260 890 404 894
rect 61 850 195 859
rect 255 850 389 859
rect 46 815 190 819
rect 46 809 190 813
rect 61 769 195 778
rect 260 815 404 819
rect 260 809 404 813
rect 46 734 190 738
rect 46 728 190 732
rect 255 769 389 778
rect 260 734 404 738
rect 260 728 404 732
rect 61 688 195 697
rect 41 653 170 657
rect 255 688 389 697
rect 280 653 409 657
<< hvpsubstratepdiff >>
rect 0 1009 450 1010
rect 0 1007 12 1009
rect 0 628 1 1007
rect 10 1000 12 1007
rect 171 1000 279 1009
rect 438 1007 450 1009
rect 438 1000 440 1007
rect 10 999 440 1000
rect 10 631 11 999
rect 439 631 440 999
rect 10 628 14 631
rect 0 627 14 628
rect 273 627 282 631
rect 436 628 440 631
rect 449 628 450 1007
rect 436 627 450 628
rect 0 620 450 627
rect 0 616 3 620
rect 447 616 450 620
rect 0 610 450 616
rect 0 606 3 610
rect 447 606 450 610
rect 0 600 450 606
rect 0 596 3 600
rect 447 596 450 600
rect 0 590 450 596
rect 0 586 3 590
rect 447 586 450 590
rect 0 580 450 586
rect 0 576 3 580
rect 447 576 450 580
rect 0 570 450 576
rect 0 566 3 570
rect 447 566 450 570
rect 0 560 450 566
rect 0 556 3 560
rect 447 556 450 560
rect 0 550 450 556
rect 0 546 3 550
rect 447 546 450 550
rect 0 540 450 546
rect 0 536 3 540
rect 447 536 450 540
rect 0 530 450 536
rect 0 526 3 530
rect 447 526 450 530
rect 0 520 450 526
rect 20 372 430 373
rect 20 363 21 372
rect 425 363 430 372
rect 20 361 430 363
rect 20 357 21 361
rect 20 351 430 357
rect 20 347 21 351
rect 20 341 430 347
rect 20 337 21 341
rect 20 331 430 337
rect 20 327 21 331
rect 20 321 430 327
rect 20 317 21 321
rect 20 311 430 317
rect 20 307 21 311
rect 20 301 430 307
rect 20 297 21 301
rect 20 291 430 297
rect 20 287 21 291
rect 20 281 430 287
rect 20 277 21 281
rect 20 271 430 277
rect 20 267 21 271
rect 20 261 430 267
rect 20 257 21 261
rect 20 251 430 257
rect 20 247 21 251
rect 20 241 430 247
rect 20 237 21 241
rect 20 231 430 237
rect 20 227 21 231
rect 20 221 430 227
rect 20 217 21 221
rect 20 211 430 217
rect 20 207 21 211
rect 20 201 430 207
rect 20 197 21 201
rect 20 191 430 197
rect 20 187 21 191
rect 20 181 430 187
rect 20 177 21 181
rect 20 171 430 177
rect 20 167 21 171
rect 20 161 430 167
rect 20 157 21 161
rect 20 151 430 157
rect 20 147 21 151
rect 20 141 430 147
rect 20 137 21 141
rect 20 131 430 137
rect 20 127 21 131
rect 20 121 430 127
rect 20 117 21 121
rect 20 111 430 117
rect 20 107 21 111
rect 20 101 430 107
rect 20 97 21 101
rect 20 91 430 97
rect 20 87 21 91
rect 20 81 430 87
rect 20 77 21 81
rect 20 71 430 77
rect 20 67 21 71
rect 20 61 430 67
rect 20 57 21 61
rect 20 51 430 57
rect 20 47 21 51
rect 20 41 430 47
rect 20 37 21 41
rect 20 31 430 37
rect 20 27 21 31
rect 20 17 430 27
<< hvnsubstratendiff >>
rect 20 988 430 990
rect 24 987 425 988
rect 24 983 40 987
rect 174 983 276 987
rect 410 983 425 987
rect 24 979 425 983
rect 24 654 30 979
rect 38 977 213 979
rect 218 925 232 979
rect 237 977 412 979
rect 218 921 223 925
rect 227 921 232 925
rect 218 915 232 921
rect 218 906 223 915
rect 227 906 232 915
rect 218 900 232 906
rect 218 891 223 900
rect 227 891 232 900
rect 218 885 232 891
rect 218 876 223 885
rect 227 876 232 885
rect 218 870 232 876
rect 218 866 223 870
rect 227 866 232 870
rect 218 834 232 866
rect 218 830 223 834
rect 227 830 232 834
rect 218 824 232 830
rect 218 815 223 824
rect 227 815 232 824
rect 218 809 232 815
rect 218 800 223 809
rect 227 800 232 809
rect 218 794 232 800
rect 218 785 223 794
rect 227 785 232 794
rect 218 779 232 785
rect 218 775 223 779
rect 227 775 232 779
rect 218 727 232 775
rect 218 723 223 727
rect 227 723 232 727
rect 218 717 232 723
rect 218 708 223 717
rect 227 708 232 717
rect 218 702 232 708
rect 218 693 223 702
rect 227 693 232 702
rect 218 687 232 693
rect 218 678 223 687
rect 227 678 232 687
rect 218 672 232 678
rect 218 668 223 672
rect 227 668 232 672
rect 20 651 30 654
rect 38 651 213 652
rect 20 642 21 651
rect 170 650 213 651
rect 218 650 232 668
rect 237 651 412 652
rect 420 654 425 979
rect 429 654 430 988
rect 420 651 430 654
rect 237 650 280 651
rect 170 642 280 650
rect 429 642 430 651
rect 20 640 430 642
rect 0 485 450 490
rect 0 484 218 485
rect 0 480 2 484
rect 131 481 218 484
rect 232 484 450 485
rect 232 481 324 484
rect 131 480 324 481
rect 448 480 450 484
rect 0 475 450 480
rect 0 474 218 475
rect 0 470 2 474
rect 131 471 218 474
rect 232 474 450 475
rect 232 471 324 474
rect 131 470 324 471
rect 448 470 450 474
rect 0 465 450 470
rect 0 464 218 465
rect 0 460 2 464
rect 131 461 218 464
rect 232 464 450 465
rect 232 461 324 464
rect 131 460 324 461
rect 448 460 450 464
rect 0 455 450 460
rect 0 454 218 455
rect 0 450 2 454
rect 131 450 218 454
rect 0 444 218 450
rect 0 440 2 444
rect 131 440 218 444
rect 0 434 218 440
rect 0 430 2 434
rect 131 430 218 434
rect 0 424 218 430
rect 0 420 2 424
rect 131 421 218 424
rect 232 454 450 455
rect 232 450 324 454
rect 448 450 450 454
rect 232 444 450 450
rect 232 440 324 444
rect 448 440 450 444
rect 232 434 450 440
rect 232 430 324 434
rect 448 430 450 434
rect 232 424 450 430
rect 232 421 324 424
rect 131 420 324 421
rect 448 420 450 424
rect 0 415 450 420
rect 0 414 218 415
rect 0 410 2 414
rect 131 411 218 414
rect 232 414 450 415
rect 232 411 324 414
rect 131 410 324 411
rect 448 410 450 414
rect 0 405 450 410
rect 0 404 218 405
rect 0 400 2 404
rect 131 401 218 404
rect 232 404 450 405
rect 232 401 324 404
rect 131 400 324 401
rect 448 400 450 404
rect 0 395 450 400
rect 0 394 218 395
rect 0 390 2 394
rect 131 391 218 394
rect 232 394 450 395
rect 232 391 324 394
rect 131 390 324 391
rect 448 390 450 394
rect 0 383 450 390
rect 0 379 12 383
rect 131 379 320 383
rect 434 379 450 383
rect 0 0 2 379
rect 11 11 13 379
rect 436 11 439 379
rect 11 9 439 11
rect 11 0 15 9
rect 169 0 281 9
rect 435 0 439 9
rect 448 0 450 379
<< hvpsubstratepcontact >>
rect 1 628 10 1007
rect 12 1000 171 1009
rect 279 1000 438 1009
rect 14 627 273 631
rect 282 627 436 631
rect 440 628 449 1007
rect 3 616 447 620
rect 3 606 447 610
rect 3 596 447 600
rect 3 586 447 590
rect 3 576 447 580
rect 3 566 447 570
rect 3 556 447 560
rect 3 546 447 550
rect 3 536 447 540
rect 3 526 447 530
rect 21 363 425 372
rect 21 357 430 361
rect 21 347 430 351
rect 21 337 430 341
rect 21 327 430 331
rect 21 317 430 321
rect 21 307 430 311
rect 21 297 430 301
rect 21 287 430 291
rect 21 277 430 281
rect 21 267 430 271
rect 21 257 430 261
rect 21 247 430 251
rect 21 237 430 241
rect 21 227 430 231
rect 21 217 430 221
rect 21 207 430 211
rect 21 197 430 201
rect 21 187 430 191
rect 21 177 430 181
rect 21 167 430 171
rect 21 157 430 161
rect 21 147 430 151
rect 21 137 430 141
rect 21 127 430 131
rect 21 117 430 121
rect 21 107 430 111
rect 21 97 430 101
rect 21 87 430 91
rect 21 77 430 81
rect 21 67 430 71
rect 21 57 430 61
rect 21 47 430 51
rect 21 37 430 41
rect 21 27 430 31
<< hvnsubstratencontact >>
rect 20 654 24 988
rect 40 983 174 987
rect 276 983 410 987
rect 223 921 227 925
rect 223 906 227 915
rect 223 891 227 900
rect 223 876 227 885
rect 223 866 227 870
rect 223 830 227 834
rect 223 815 227 824
rect 223 800 227 809
rect 223 785 227 794
rect 223 775 227 779
rect 223 723 227 727
rect 223 708 227 717
rect 223 693 227 702
rect 223 678 227 687
rect 223 668 227 672
rect 21 642 170 651
rect 425 654 429 988
rect 280 642 429 651
rect 2 480 131 484
rect 218 481 232 485
rect 324 480 448 484
rect 2 470 131 474
rect 218 471 232 475
rect 324 470 448 474
rect 2 460 131 464
rect 218 461 232 465
rect 324 460 448 464
rect 2 450 131 454
rect 2 440 131 444
rect 2 430 131 434
rect 2 420 131 424
rect 218 421 232 455
rect 324 450 448 454
rect 324 440 448 444
rect 324 430 448 434
rect 324 420 448 424
rect 2 410 131 414
rect 218 411 232 415
rect 324 410 448 414
rect 2 400 131 404
rect 218 401 232 405
rect 324 400 448 404
rect 2 390 131 394
rect 218 391 232 395
rect 324 390 448 394
rect 12 379 131 383
rect 320 379 434 383
rect 2 0 11 379
rect 15 0 169 9
rect 281 0 435 9
rect 439 0 448 379
<< polysilicon >>
rect 31 966 38 968
rect 31 662 32 966
rect 36 965 38 966
rect 213 965 216 968
rect 36 907 37 965
rect 234 965 237 968
rect 412 966 419 968
rect 412 965 414 966
rect 36 904 38 907
rect 213 904 216 907
rect 413 907 414 965
rect 36 886 37 904
rect 234 904 237 907
rect 412 904 414 907
rect 36 883 38 886
rect 213 883 216 886
rect 413 886 414 904
rect 36 826 37 883
rect 234 883 237 886
rect 412 883 414 886
rect 36 823 38 826
rect 213 823 216 826
rect 413 826 414 883
rect 36 805 37 823
rect 234 823 237 826
rect 412 823 414 826
rect 36 802 38 805
rect 213 802 216 805
rect 36 745 37 802
rect 413 805 414 823
rect 234 802 237 805
rect 412 802 414 805
rect 36 742 38 745
rect 213 742 216 745
rect 36 724 37 742
rect 413 745 414 802
rect 234 742 237 745
rect 412 742 414 745
rect 36 721 38 724
rect 213 721 216 724
rect 413 724 414 742
rect 36 664 37 721
rect 234 721 237 724
rect 412 721 414 724
rect 36 662 38 664
rect 31 661 38 662
rect 213 661 216 664
rect 413 664 414 721
rect 234 661 237 664
rect 412 662 414 664
rect 418 662 419 966
rect 412 661 419 662
<< polycontact >>
rect 32 662 36 966
rect 414 662 418 966
<< metal1 >>
rect 30 1495 420 1500
rect 30 1114 34 1495
rect 415 1114 420 1495
rect 30 1110 420 1114
rect 137 1100 313 1110
rect 147 1090 303 1100
rect 157 1080 293 1090
rect 167 1070 283 1080
rect 0 1009 174 1010
rect 0 1007 12 1009
rect 0 628 1 1007
rect 10 1000 12 1007
rect 171 1000 174 1009
rect 10 999 174 1000
rect 10 631 11 999
rect 178 998 272 1070
rect 276 1009 450 1010
rect 276 1000 279 1009
rect 438 1007 450 1009
rect 438 1000 440 1007
rect 276 999 440 1000
rect 20 988 174 989
rect 24 654 25 988
rect 29 987 174 988
rect 29 983 40 987
rect 181 984 269 998
rect 276 988 430 989
rect 276 987 420 988
rect 29 982 174 983
rect 29 978 40 982
rect 29 976 174 978
rect 29 972 41 976
rect 170 972 174 976
rect 29 966 174 972
rect 186 969 264 984
rect 410 983 420 987
rect 276 982 420 983
rect 410 978 420 982
rect 276 976 420 978
rect 276 972 280 976
rect 409 972 420 976
rect 29 662 32 966
rect 36 964 174 966
rect 36 940 39 964
rect 48 960 52 964
rect 166 960 174 964
rect 48 940 51 960
rect 199 957 251 969
rect 276 966 420 972
rect 276 964 414 966
rect 276 960 284 964
rect 398 960 402 964
rect 36 938 51 940
rect 36 934 39 938
rect 48 934 51 938
rect 36 932 51 934
rect 36 908 39 932
rect 48 912 51 932
rect 56 941 394 957
rect 56 937 61 941
rect 195 937 255 941
rect 389 937 394 941
rect 56 935 394 937
rect 56 931 61 935
rect 195 931 255 935
rect 389 931 394 935
rect 56 928 394 931
rect 56 915 220 928
rect 48 908 52 912
rect 186 908 195 912
rect 36 900 195 908
rect 36 896 46 900
rect 190 896 195 900
rect 36 894 195 896
rect 36 890 46 894
rect 190 890 195 894
rect 36 882 195 890
rect 36 853 39 882
rect 48 878 52 882
rect 186 878 195 882
rect 48 853 51 878
rect 199 875 220 915
rect 36 851 51 853
rect 36 827 39 851
rect 48 831 51 851
rect 56 863 220 875
rect 223 920 227 921
rect 223 915 227 916
rect 223 905 227 906
rect 223 900 227 901
rect 223 890 227 891
rect 223 885 227 886
rect 223 875 227 876
rect 223 870 227 871
rect 230 915 394 928
rect 399 940 402 960
rect 411 940 414 964
rect 399 938 414 940
rect 399 934 402 938
rect 411 934 414 938
rect 399 932 414 934
rect 230 875 251 915
rect 399 912 402 932
rect 255 908 264 912
rect 398 908 402 912
rect 411 908 414 932
rect 255 900 414 908
rect 255 896 260 900
rect 404 896 414 900
rect 255 894 414 896
rect 255 890 260 894
rect 404 890 414 894
rect 255 882 414 890
rect 255 878 264 882
rect 398 878 402 882
rect 230 863 394 875
rect 56 859 394 863
rect 56 850 61 859
rect 195 850 255 859
rect 389 850 394 859
rect 56 837 394 850
rect 56 834 220 837
rect 230 834 394 837
rect 399 853 402 878
rect 411 853 414 882
rect 399 851 414 853
rect 48 827 52 831
rect 186 827 195 831
rect 36 819 195 827
rect 36 815 46 819
rect 190 815 195 819
rect 36 813 195 815
rect 36 809 46 813
rect 190 809 195 813
rect 36 801 195 809
rect 36 772 39 801
rect 48 797 52 801
rect 186 797 195 801
rect 48 772 51 797
rect 199 794 220 834
rect 36 770 51 772
rect 36 746 39 770
rect 48 750 51 770
rect 56 778 220 794
rect 56 769 61 778
rect 195 772 220 778
rect 223 829 227 830
rect 223 824 227 825
rect 223 814 227 815
rect 223 809 227 810
rect 223 799 227 800
rect 223 794 227 795
rect 223 784 227 785
rect 223 779 227 780
rect 230 794 251 834
rect 399 831 402 851
rect 255 827 264 831
rect 398 827 402 831
rect 411 827 414 851
rect 255 819 414 827
rect 255 815 260 819
rect 404 815 414 819
rect 255 813 414 815
rect 255 809 260 813
rect 404 809 414 813
rect 255 801 414 809
rect 255 797 264 801
rect 398 797 402 801
rect 230 778 394 794
rect 230 772 255 778
rect 195 769 255 772
rect 389 769 394 778
rect 56 753 394 769
rect 399 772 402 797
rect 411 772 414 801
rect 399 770 414 772
rect 48 746 52 750
rect 186 746 195 750
rect 36 738 195 746
rect 36 734 46 738
rect 190 734 195 738
rect 36 732 195 734
rect 36 728 46 732
rect 190 728 195 732
rect 36 720 195 728
rect 36 691 39 720
rect 48 716 52 720
rect 186 716 195 720
rect 199 730 251 753
rect 399 750 402 770
rect 48 691 51 716
rect 199 713 220 730
rect 36 689 51 691
rect 36 665 39 689
rect 48 669 51 689
rect 56 697 220 713
rect 56 688 61 697
rect 195 688 220 697
rect 56 672 220 688
rect 48 665 52 669
rect 166 665 174 669
rect 36 662 174 665
rect 29 657 174 662
rect 29 654 41 657
rect 20 653 41 654
rect 170 653 174 657
rect 20 651 174 653
rect 20 642 21 651
rect 170 642 174 651
rect 20 641 174 642
rect 178 665 220 672
rect 223 722 227 723
rect 223 717 227 718
rect 223 707 227 708
rect 223 702 227 703
rect 223 692 227 693
rect 223 687 227 688
rect 223 677 227 678
rect 223 672 227 673
rect 230 713 251 730
rect 255 746 264 750
rect 398 746 402 750
rect 411 746 414 770
rect 255 738 414 746
rect 255 734 260 738
rect 404 734 414 738
rect 255 732 414 734
rect 255 728 260 732
rect 404 728 414 732
rect 255 720 414 728
rect 255 716 264 720
rect 398 716 402 720
rect 230 697 394 713
rect 230 688 255 697
rect 389 688 394 697
rect 230 672 394 688
rect 399 691 402 716
rect 411 691 414 720
rect 399 689 414 691
rect 230 665 272 672
rect 399 669 402 689
rect 178 631 272 665
rect 276 665 284 669
rect 398 665 402 669
rect 411 665 414 689
rect 276 662 414 665
rect 418 662 420 966
rect 276 657 420 662
rect 276 653 280 657
rect 409 654 420 657
rect 424 654 425 988
rect 429 654 430 988
rect 409 653 430 654
rect 276 651 430 653
rect 276 642 280 651
rect 429 642 430 651
rect 276 641 430 642
rect 439 631 440 999
rect 10 628 14 631
rect 0 627 14 628
rect 273 627 282 631
rect 436 628 440 631
rect 449 628 450 1007
rect 436 627 450 628
rect 0 625 450 627
rect 0 621 3 625
rect 447 621 450 625
rect 0 620 450 621
rect 0 616 3 620
rect 447 616 450 620
rect 0 615 450 616
rect 0 611 3 615
rect 447 611 450 615
rect 0 610 450 611
rect 0 606 3 610
rect 447 606 450 610
rect 0 605 450 606
rect 0 601 3 605
rect 447 601 450 605
rect 0 600 450 601
rect 0 596 3 600
rect 447 596 450 600
rect 0 595 450 596
rect 0 591 3 595
rect 447 591 450 595
rect 0 590 450 591
rect 0 586 3 590
rect 447 586 450 590
rect 0 585 450 586
rect 0 581 3 585
rect 447 581 450 585
rect 0 580 450 581
rect 0 576 3 580
rect 447 576 450 580
rect 0 575 450 576
rect 0 571 3 575
rect 447 571 450 575
rect 0 570 450 571
rect 0 566 3 570
rect 447 566 450 570
rect 0 565 450 566
rect 0 561 3 565
rect 447 561 450 565
rect 0 560 450 561
rect 0 556 3 560
rect 447 556 450 560
rect 0 555 450 556
rect 0 551 3 555
rect 447 551 450 555
rect 0 550 450 551
rect 0 546 3 550
rect 447 546 450 550
rect 0 545 450 546
rect 0 541 3 545
rect 447 541 450 545
rect 0 540 450 541
rect 0 536 3 540
rect 447 536 450 540
rect 0 535 450 536
rect 0 531 3 535
rect 447 531 450 535
rect 0 530 450 531
rect 0 526 3 530
rect 447 526 450 530
rect 0 525 450 526
rect 0 521 3 525
rect 447 521 450 525
rect 0 485 2 489
rect 0 484 131 485
rect 0 480 2 484
rect 0 479 131 480
rect 0 475 2 479
rect 0 474 131 475
rect 0 470 2 474
rect 0 469 131 470
rect 0 465 2 469
rect 0 464 131 465
rect 0 460 2 464
rect 0 459 131 460
rect 0 455 2 459
rect 0 454 131 455
rect 0 450 2 454
rect 0 449 131 450
rect 0 445 2 449
rect 0 444 131 445
rect 0 440 2 444
rect 0 439 131 440
rect 0 435 2 439
rect 0 434 131 435
rect 0 430 2 434
rect 0 429 131 430
rect 0 425 2 429
rect 0 424 131 425
rect 0 420 2 424
rect 0 419 131 420
rect 0 415 2 419
rect 0 414 131 415
rect 0 410 2 414
rect 0 409 131 410
rect 0 405 2 409
rect 0 404 131 405
rect 0 400 2 404
rect 0 399 131 400
rect 0 395 2 399
rect 0 394 131 395
rect 0 390 2 394
rect 0 389 131 390
rect 0 385 2 389
rect 0 383 131 385
rect 0 379 12 383
rect 0 0 2 379
rect 11 11 13 379
rect 135 372 173 521
rect 177 372 215 521
rect 218 485 232 486
rect 218 480 232 481
rect 218 475 232 476
rect 218 470 232 471
rect 218 465 232 466
rect 218 460 232 461
rect 218 455 232 456
rect 218 420 232 421
rect 218 415 232 416
rect 218 410 232 411
rect 218 405 232 406
rect 218 400 232 401
rect 218 395 232 396
rect 218 390 232 391
rect 236 372 274 521
rect 278 372 316 521
rect 320 485 324 489
rect 448 485 450 489
rect 320 484 450 485
rect 320 480 324 484
rect 448 480 450 484
rect 320 479 450 480
rect 320 475 324 479
rect 448 475 450 479
rect 320 474 450 475
rect 320 470 324 474
rect 448 470 450 474
rect 320 469 450 470
rect 320 465 324 469
rect 448 465 450 469
rect 320 464 450 465
rect 320 460 324 464
rect 448 460 450 464
rect 320 459 450 460
rect 320 455 324 459
rect 448 455 450 459
rect 320 454 450 455
rect 320 450 324 454
rect 448 450 450 454
rect 320 449 450 450
rect 320 445 324 449
rect 448 445 450 449
rect 320 444 450 445
rect 320 440 324 444
rect 448 440 450 444
rect 320 439 450 440
rect 320 435 324 439
rect 448 435 450 439
rect 320 434 450 435
rect 320 430 324 434
rect 448 430 450 434
rect 320 429 450 430
rect 320 425 324 429
rect 448 425 450 429
rect 320 424 450 425
rect 320 420 324 424
rect 448 420 450 424
rect 320 419 450 420
rect 320 415 324 419
rect 448 415 450 419
rect 320 414 450 415
rect 320 410 324 414
rect 448 410 450 414
rect 320 409 450 410
rect 320 405 324 409
rect 448 405 450 409
rect 320 404 450 405
rect 320 400 324 404
rect 448 400 450 404
rect 320 399 450 400
rect 320 395 324 399
rect 448 395 450 399
rect 320 394 450 395
rect 320 390 324 394
rect 448 390 450 394
rect 320 389 450 390
rect 320 385 324 389
rect 448 385 450 389
rect 320 383 450 385
rect 434 379 450 383
rect 425 363 429 372
rect 21 361 429 363
rect 21 356 430 357
rect 21 351 430 352
rect 21 346 430 347
rect 21 341 430 342
rect 21 336 430 337
rect 21 331 430 332
rect 21 326 430 327
rect 21 321 430 322
rect 21 316 430 317
rect 21 311 430 312
rect 21 306 430 307
rect 21 301 430 302
rect 21 296 430 297
rect 21 291 430 292
rect 21 286 430 287
rect 21 281 430 282
rect 21 276 430 277
rect 21 271 430 272
rect 21 266 430 267
rect 21 261 430 262
rect 21 256 430 257
rect 21 251 430 252
rect 21 246 430 247
rect 21 241 430 242
rect 21 236 430 237
rect 21 231 430 232
rect 21 226 430 227
rect 21 221 430 222
rect 21 216 430 217
rect 21 211 430 212
rect 21 206 430 207
rect 21 201 430 202
rect 21 196 430 197
rect 21 191 430 192
rect 21 186 430 187
rect 21 181 430 182
rect 21 176 430 177
rect 21 171 430 172
rect 21 166 430 167
rect 21 161 430 162
rect 21 156 430 157
rect 21 151 430 152
rect 21 146 430 147
rect 21 141 430 142
rect 21 136 430 137
rect 21 131 430 132
rect 21 126 430 127
rect 21 121 430 122
rect 21 116 430 117
rect 21 111 430 112
rect 21 106 430 107
rect 21 101 430 102
rect 21 96 430 97
rect 21 91 430 92
rect 21 86 430 87
rect 21 81 430 82
rect 21 76 430 77
rect 21 71 430 72
rect 21 66 430 67
rect 21 61 430 62
rect 21 56 430 57
rect 21 51 430 52
rect 21 46 430 47
rect 21 41 430 42
rect 21 36 430 37
rect 21 31 430 32
rect 21 26 430 27
rect 21 18 429 22
rect 11 9 171 11
rect 11 0 15 9
rect 169 0 171 9
rect 174 0 274 18
rect 436 11 439 379
rect 278 9 439 11
rect 278 0 281 9
rect 435 0 439 9
rect 448 0 450 379
<< m2contact >>
rect 25 654 29 988
rect 40 978 174 982
rect 276 978 410 982
rect 39 940 48 964
rect 52 960 166 964
rect 284 960 398 964
rect 39 934 48 938
rect 39 908 48 932
rect 52 908 186 912
rect 39 853 48 882
rect 52 878 186 882
rect 39 827 48 851
rect 223 916 227 920
rect 223 901 227 905
rect 223 886 227 890
rect 223 871 227 875
rect 402 940 411 964
rect 402 934 411 938
rect 264 908 398 912
rect 402 908 411 932
rect 264 878 398 882
rect 402 853 411 882
rect 52 827 186 831
rect 39 772 48 801
rect 52 797 186 801
rect 39 746 48 770
rect 223 825 227 829
rect 223 810 227 814
rect 223 795 227 799
rect 223 780 227 784
rect 264 827 398 831
rect 402 827 411 851
rect 264 797 398 801
rect 402 772 411 801
rect 52 746 186 750
rect 39 691 48 720
rect 52 716 186 720
rect 39 665 48 689
rect 52 665 166 669
rect 223 718 227 722
rect 223 703 227 707
rect 223 688 227 692
rect 223 673 227 677
rect 264 746 398 750
rect 402 746 411 770
rect 264 716 398 720
rect 402 691 411 720
rect 284 665 398 669
rect 402 665 411 689
rect 420 654 424 988
rect 3 621 447 625
rect 3 611 447 615
rect 3 601 447 605
rect 3 591 447 595
rect 3 581 447 585
rect 3 571 447 575
rect 3 561 447 565
rect 3 551 447 555
rect 3 541 447 545
rect 3 531 447 535
rect 3 521 447 525
rect 2 485 131 489
rect 2 475 131 479
rect 2 465 131 469
rect 2 455 131 459
rect 2 445 131 449
rect 2 435 131 439
rect 2 425 131 429
rect 2 415 131 419
rect 2 405 131 409
rect 2 395 131 399
rect 2 385 131 389
rect 218 476 232 480
rect 218 466 232 470
rect 218 456 232 460
rect 218 416 232 420
rect 218 406 232 410
rect 218 396 232 400
rect 324 485 448 489
rect 324 475 448 479
rect 324 465 448 469
rect 324 455 448 459
rect 324 445 448 449
rect 324 435 448 439
rect 324 425 448 429
rect 324 415 448 419
rect 324 405 448 409
rect 324 395 448 399
rect 324 385 448 389
rect 21 352 430 356
rect 21 342 430 346
rect 21 332 430 336
rect 21 322 430 326
rect 21 312 430 316
rect 21 302 430 306
rect 21 292 430 296
rect 21 282 430 286
rect 21 272 430 276
rect 21 262 430 266
rect 21 252 430 256
rect 21 242 430 246
rect 21 232 430 236
rect 21 222 430 226
rect 21 212 430 216
rect 21 202 430 206
rect 21 192 430 196
rect 21 182 430 186
rect 21 172 430 176
rect 21 162 430 166
rect 21 152 430 156
rect 21 142 430 146
rect 21 132 430 136
rect 21 122 430 126
rect 21 112 430 116
rect 21 102 430 106
rect 21 92 430 96
rect 21 82 430 86
rect 21 72 430 76
rect 21 62 430 66
rect 21 52 430 56
rect 21 42 430 46
rect 21 32 430 36
rect 21 22 430 26
<< metal2 >>
rect 30 1495 420 1500
rect 30 1114 34 1495
rect 415 1114 420 1495
rect 30 1110 420 1114
rect 0 988 450 1010
rect 0 654 25 988
rect 29 982 420 988
rect 29 978 40 982
rect 174 978 276 982
rect 410 978 420 982
rect 29 964 420 978
rect 29 940 39 964
rect 48 960 52 964
rect 166 960 284 964
rect 398 960 402 964
rect 48 940 402 960
rect 411 940 420 964
rect 29 938 420 940
rect 29 934 39 938
rect 48 934 402 938
rect 411 934 420 938
rect 29 932 420 934
rect 29 908 39 932
rect 48 920 402 932
rect 48 916 223 920
rect 227 916 402 920
rect 48 912 402 916
rect 48 908 52 912
rect 186 908 264 912
rect 398 908 402 912
rect 411 908 420 932
rect 29 905 420 908
rect 29 901 223 905
rect 227 901 420 905
rect 29 890 420 901
rect 29 886 223 890
rect 227 886 420 890
rect 29 882 420 886
rect 29 853 39 882
rect 48 878 52 882
rect 186 878 264 882
rect 398 878 402 882
rect 48 875 402 878
rect 48 871 223 875
rect 227 871 402 875
rect 48 853 402 871
rect 411 853 420 882
rect 29 851 420 853
rect 29 827 39 851
rect 48 831 402 851
rect 48 827 52 831
rect 186 829 264 831
rect 186 827 223 829
rect 29 825 223 827
rect 227 827 264 829
rect 398 827 402 831
rect 411 827 420 851
rect 227 825 420 827
rect 29 814 420 825
rect 29 810 223 814
rect 227 810 420 814
rect 29 801 420 810
rect 29 772 39 801
rect 48 797 52 801
rect 186 799 264 801
rect 186 797 223 799
rect 48 795 223 797
rect 227 797 264 799
rect 398 797 402 801
rect 227 795 402 797
rect 48 784 402 795
rect 48 780 223 784
rect 227 780 402 784
rect 48 772 402 780
rect 411 772 420 801
rect 29 770 420 772
rect 29 746 39 770
rect 48 750 402 770
rect 48 746 52 750
rect 186 746 264 750
rect 398 746 402 750
rect 411 746 420 770
rect 29 722 420 746
rect 29 720 223 722
rect 29 691 39 720
rect 48 716 52 720
rect 186 718 223 720
rect 227 720 420 722
rect 227 718 264 720
rect 186 716 264 718
rect 398 716 402 720
rect 48 707 402 716
rect 48 703 223 707
rect 227 703 402 707
rect 48 692 402 703
rect 48 691 223 692
rect 29 689 223 691
rect 29 665 39 689
rect 48 688 223 689
rect 227 691 402 692
rect 411 691 420 720
rect 227 689 420 691
rect 227 688 402 689
rect 48 677 402 688
rect 48 673 223 677
rect 227 673 402 677
rect 48 669 402 673
rect 48 665 52 669
rect 166 665 284 669
rect 398 665 402 669
rect 411 665 420 689
rect 29 654 420 665
rect 424 654 450 988
rect 0 648 450 654
rect 0 625 450 626
rect 0 621 3 625
rect 447 621 450 625
rect 0 615 450 621
rect 0 611 3 615
rect 447 611 450 615
rect 0 605 450 611
rect 0 601 3 605
rect 447 601 450 605
rect 0 595 450 601
rect 0 591 3 595
rect 447 591 450 595
rect 0 585 450 591
rect 0 581 3 585
rect 447 581 450 585
rect 0 575 450 581
rect 0 571 3 575
rect 447 571 450 575
rect 0 565 450 571
rect 0 561 3 565
rect 447 561 450 565
rect 0 555 450 561
rect 0 551 3 555
rect 447 551 450 555
rect 0 545 450 551
rect 0 541 3 545
rect 447 541 450 545
rect 0 535 450 541
rect 0 531 3 535
rect 447 531 450 535
rect 0 525 450 531
rect 0 521 3 525
rect 447 521 450 525
rect 0 485 2 489
rect 131 485 324 489
rect 448 485 450 489
rect 0 480 450 485
rect 0 479 218 480
rect 0 475 2 479
rect 131 476 218 479
rect 232 479 450 480
rect 232 476 324 479
rect 131 475 324 476
rect 448 475 450 479
rect 0 470 450 475
rect 0 469 218 470
rect 0 465 2 469
rect 131 466 218 469
rect 232 469 450 470
rect 232 466 324 469
rect 131 465 324 466
rect 448 465 450 469
rect 0 460 450 465
rect 0 459 218 460
rect 0 455 2 459
rect 131 456 218 459
rect 232 459 450 460
rect 232 456 324 459
rect 131 455 324 456
rect 448 455 450 459
rect 0 449 450 455
rect 0 445 2 449
rect 131 445 324 449
rect 448 445 450 449
rect 0 439 450 445
rect 0 435 2 439
rect 131 435 324 439
rect 448 435 450 439
rect 0 429 450 435
rect 0 425 2 429
rect 131 425 324 429
rect 448 425 450 429
rect 0 420 450 425
rect 0 419 218 420
rect 0 415 2 419
rect 131 416 218 419
rect 232 419 450 420
rect 232 416 324 419
rect 131 415 324 416
rect 448 415 450 419
rect 0 410 450 415
rect 0 409 218 410
rect 0 405 2 409
rect 131 406 218 409
rect 232 409 450 410
rect 232 406 324 409
rect 131 405 324 406
rect 448 405 450 409
rect 0 400 450 405
rect 0 399 218 400
rect 0 395 2 399
rect 131 396 218 399
rect 232 399 450 400
rect 232 396 324 399
rect 131 395 324 396
rect 448 395 450 399
rect 0 389 450 395
rect 0 385 2 389
rect 131 385 324 389
rect 448 385 450 389
rect 0 384 450 385
rect 440 383 448 384
rect 0 356 450 362
rect 0 352 21 356
rect 430 352 450 356
rect 0 346 450 352
rect 0 342 21 346
rect 430 342 450 346
rect 0 336 450 342
rect 0 332 21 336
rect 430 332 450 336
rect 0 326 450 332
rect 0 322 21 326
rect 430 322 450 326
rect 0 316 450 322
rect 0 312 21 316
rect 430 312 450 316
rect 0 306 450 312
rect 0 302 21 306
rect 430 302 450 306
rect 0 296 450 302
rect 0 292 21 296
rect 430 292 450 296
rect 0 286 450 292
rect 0 282 21 286
rect 430 282 450 286
rect 0 276 450 282
rect 0 272 21 276
rect 430 272 450 276
rect 0 266 450 272
rect 0 262 21 266
rect 430 262 450 266
rect 0 256 450 262
rect 0 252 21 256
rect 430 252 450 256
rect 0 246 450 252
rect 0 242 21 246
rect 430 242 450 246
rect 0 236 450 242
rect 0 232 21 236
rect 430 232 450 236
rect 0 226 450 232
rect 0 222 21 226
rect 430 222 450 226
rect 0 216 450 222
rect 0 212 21 216
rect 430 212 450 216
rect 0 206 450 212
rect 0 202 21 206
rect 430 202 450 206
rect 0 196 450 202
rect 0 192 21 196
rect 430 192 450 196
rect 0 186 450 192
rect 0 182 21 186
rect 430 182 450 186
rect 0 176 450 182
rect 0 172 21 176
rect 430 172 450 176
rect 0 166 450 172
rect 0 162 21 166
rect 430 162 450 166
rect 0 156 450 162
rect 0 152 21 156
rect 430 152 450 156
rect 0 146 450 152
rect 0 142 21 146
rect 430 142 450 146
rect 0 136 450 142
rect 0 132 21 136
rect 430 132 450 136
rect 0 126 450 132
rect 0 122 21 126
rect 430 122 450 126
rect 0 116 450 122
rect 0 112 21 116
rect 430 112 450 116
rect 0 106 450 112
rect 0 102 21 106
rect 430 102 450 106
rect 0 96 450 102
rect 0 92 21 96
rect 430 92 450 96
rect 0 86 450 92
rect 0 82 21 86
rect 430 82 450 86
rect 0 76 450 82
rect 0 72 21 76
rect 430 72 450 76
rect 0 66 450 72
rect 0 62 21 66
rect 430 62 450 66
rect 0 56 450 62
rect 0 52 21 56
rect 430 52 450 56
rect 0 46 450 52
rect 0 42 21 46
rect 430 42 450 46
rect 0 36 450 42
rect 0 32 21 36
rect 430 32 450 36
rect 0 26 450 32
rect 0 22 21 26
rect 430 22 450 26
rect 0 0 450 22
<< pad >>
rect 34 1114 415 1495
<< m1p >>
rect 174 0 274 4
<< m4p >>
rect 187 1274 256 1349
<< labels >>
rlabel metal1 224 0 224 0 8 gnd
rlabel m4p 218 1310 218 1310 1 YPAD
<< end >>

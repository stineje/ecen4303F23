magic
tech sky130A
magscale 1 2
timestamp 1701189950
<< nwell >>
rect 24 370 478 657
<< nmos >>
rect 124 110 154 194
rect 342 110 372 194
<< pmos >>
rect 124 406 154 490
rect 342 406 372 490
<< ndiff >>
rect 51 154 124 194
rect 51 118 76 154
rect 110 118 124 154
rect 51 110 124 118
rect 154 154 215 194
rect 154 118 165 154
rect 199 118 215 154
rect 154 110 215 118
rect 269 154 342 194
rect 269 118 294 154
rect 328 118 342 154
rect 269 110 342 118
rect 372 154 433 194
rect 372 118 383 154
rect 417 118 433 154
rect 372 110 433 118
<< pdiff >>
rect 67 482 124 490
rect 67 446 79 482
rect 113 446 124 482
rect 67 406 124 446
rect 154 482 211 490
rect 154 446 165 482
rect 199 446 211 482
rect 154 406 211 446
rect 285 482 342 490
rect 285 446 297 482
rect 331 446 342 482
rect 285 406 342 446
rect 372 482 429 490
rect 372 446 383 482
rect 417 446 429 482
rect 372 406 429 446
<< ndiffc >>
rect 76 118 110 154
rect 165 118 199 154
rect 294 118 328 154
rect 383 118 417 154
<< pdiffc >>
rect 79 446 113 482
rect 165 446 199 482
rect 297 446 331 482
rect 383 446 417 482
<< psubdiff >>
rect 107 9 131 45
rect 167 9 191 45
rect 325 9 349 45
rect 385 9 409 45
<< nsubdiff >>
rect 102 555 126 591
rect 162 555 186 591
rect 320 555 344 591
rect 380 555 404 591
<< psubdiffcont >>
rect 131 9 167 45
rect 349 9 385 45
<< nsubdiffcont >>
rect 126 555 162 591
rect 344 555 380 591
<< poly >>
rect 124 490 154 532
rect 342 490 372 532
rect 124 364 154 406
rect 342 364 372 406
rect 124 301 154 306
rect 342 301 372 306
rect 60 285 154 301
rect 60 242 76 285
rect 124 242 154 285
rect 60 226 154 242
rect 278 285 372 301
rect 278 242 294 285
rect 342 242 372 285
rect 278 226 372 242
rect 124 194 154 226
rect 342 194 372 226
rect 124 78 154 110
rect 342 78 372 110
<< polycont >>
rect 76 242 124 285
rect 294 242 342 285
<< locali >>
rect 232 603 268 604
rect 2 591 508 603
rect 2 555 126 591
rect 162 555 344 591
rect 380 555 508 591
rect 2 534 508 555
rect 79 482 113 534
rect 79 430 113 446
rect 165 482 199 499
rect 165 364 199 446
rect 297 482 331 534
rect 297 430 331 446
rect 383 482 417 499
rect 383 364 417 446
rect 165 301 199 306
rect 2 285 124 301
rect 2 242 76 285
rect 2 226 124 242
rect 165 285 342 301
rect 165 242 294 285
rect 165 226 342 242
rect 383 290 417 306
rect 383 226 508 290
rect 76 154 110 170
rect 76 61 110 118
rect 165 154 199 226
rect 165 98 199 118
rect 294 154 328 170
rect 294 61 328 118
rect 383 154 417 226
rect 383 98 417 118
rect 2 45 508 61
rect 2 9 131 45
rect 167 9 349 45
rect 385 9 508 45
rect 2 -8 508 9
<< labels >>
rlabel locali 26 262 26 262 0 A
port 1 e
rlabel locali 460 260 460 260 0 Y
port 2 w
rlabel locali 236 26 236 26 1 gnd
port 4 n
rlabel locali 404 286 404 286 1 inv_1.Y
rlabel locali 318 264 318 264 1 inv_1.A
rlabel locali 367 27 367 27 1 inv_1.GND
rlabel locali 186 286 186 286 1 inv_0.Y
rlabel locali 100 264 100 264 1 inv_0.A
rlabel locali 149 27 149 27 1 inv_0.GND
rlabel locali 244 570 244 570 0 vdd
port 3 n
rlabel nsubdiffcont 359 573 359 573 1 inv_1.VDD
rlabel nsubdiffcont 141 573 141 573 1 inv_0.VDD
<< end >>

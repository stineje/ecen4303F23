iit018_stdcells.lef

magic
tech scmos
timestamp 1091052278
<< hvnwell >>
rect 1007 -3 1503 492
<< hvpwell >>
rect 487 517 1503 1013
rect 487 -3 983 517
<< hvpsubstratepdiff >>
rect 490 1008 1500 1010
rect 490 649 491 1008
rect 1495 649 1500 1008
rect 490 627 1500 649
rect 490 3 491 627
rect 850 520 1500 627
rect 850 3 980 520
rect 490 0 980 3
<< hvnsubstratendiff >>
rect 1010 361 1500 489
rect 1010 2 1139 361
rect 1498 2 1500 361
rect 1010 0 1500 2
<< hvpsubstratepcontact >>
rect 491 649 1495 1008
rect 491 3 850 627
<< hvnsubstratencontact >>
rect 1139 2 1498 361
<< metal1 >>
rect 490 1008 1500 1010
rect 490 649 491 1008
rect 1495 649 1500 1008
rect 490 627 1500 649
rect 490 3 491 627
rect 850 624 1500 627
rect 850 520 874 624
rect 1498 520 1500 624
rect 850 514 979 520
rect 850 5 874 514
rect 978 5 979 514
rect 850 3 979 5
rect 490 0 979 3
rect 1011 488 1500 489
rect 1495 384 1500 488
rect 1011 379 1500 384
rect 1115 361 1500 379
rect 1115 5 1139 361
rect 1011 2 1139 5
rect 1498 2 1500 361
rect 1011 0 1500 2
<< m2contact >>
rect 874 520 1498 624
rect 874 5 978 514
rect 1011 384 1495 488
rect 1011 5 1115 379
<< metal2 >>
rect 490 648 1500 1010
rect 490 0 852 648
rect 874 624 1500 626
rect 1498 520 1500 624
rect 874 514 979 520
rect 978 5 979 514
rect 874 0 979 5
rect 1011 488 1500 489
rect 1495 384 1500 488
rect 1011 379 1116 384
rect 1115 5 1116 379
rect 1011 0 1116 5
rect 1138 0 1500 362
<< end >>

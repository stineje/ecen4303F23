magic
tech scmos
timestamp 1111202490
<< metal1 >>
rect 19 706 459 710
rect 26 699 452 703
rect 12 692 28 696
rect 436 654 452 658
rect 5 614 8 618
rect 12 614 27 618
rect 436 589 459 593
rect 5 564 8 568
rect 12 564 31 568
rect 436 524 452 528
rect 12 484 31 488
rect 436 459 459 463
rect 12 434 33 437
rect 437 394 452 398
rect 12 354 28 358
rect 438 329 459 333
rect 12 303 33 307
rect 438 264 452 268
rect 12 224 30 228
rect 438 199 459 203
rect 12 174 31 177
rect 444 133 452 138
rect 12 107 20 110
rect 446 81 459 86
rect 448 23 452 27
rect 26 15 452 19
rect 19 8 459 12
<< m2contact >>
rect 15 706 19 710
rect 459 706 463 710
rect 22 699 26 703
rect 452 699 456 703
rect 8 692 12 696
rect 452 654 456 658
rect 8 614 12 618
rect 459 589 463 593
rect 8 564 12 568
rect 452 524 456 528
rect 8 484 12 488
rect 459 459 463 463
rect 8 433 12 437
rect 452 394 456 398
rect 8 354 12 358
rect 459 329 463 333
rect 8 303 12 307
rect 452 264 456 268
rect 8 224 12 228
rect 459 199 463 203
rect 8 173 12 177
rect 452 133 456 138
rect 8 106 12 110
rect 459 81 463 86
rect 452 23 456 27
rect 22 15 26 19
rect 452 15 456 19
rect 15 8 19 12
rect 459 8 463 12
<< metal2 >>
rect 5 692 8 696
rect 5 614 8 618
rect 5 564 8 568
rect 5 484 8 488
rect 5 433 8 437
rect 5 354 8 358
rect 5 303 8 307
rect 5 224 8 228
rect 5 173 8 177
rect 5 106 8 110
rect 15 12 19 706
rect 5 8 15 12
rect 22 19 26 699
rect 452 658 456 699
rect 452 528 456 654
rect 452 398 456 524
rect 452 268 456 394
rect 452 138 456 264
rect 452 27 456 133
rect 22 5 26 15
rect 44 5 47 22
rect 67 5 71 18
rect 97 5 100 23
rect 120 5 124 19
rect 150 5 153 20
rect 173 5 177 20
rect 203 5 206 21
rect 226 5 230 20
rect 256 5 259 19
rect 279 5 283 20
rect 309 5 312 19
rect 332 5 336 19
rect 362 5 365 19
rect 385 5 389 20
rect 415 5 418 20
rect 438 5 442 20
rect 452 19 456 23
rect 459 593 463 706
rect 459 463 463 589
rect 459 333 463 459
rect 459 203 463 329
rect 459 86 463 199
rect 459 12 463 81
<< m3contact >>
rect 1 692 5 696
rect 1 614 5 618
rect 1 564 5 568
rect 1 484 5 488
rect 1 433 5 437
rect 1 354 5 358
rect 1 303 5 307
rect 1 224 5 228
rect 1 173 5 177
rect 1 106 5 110
rect 1 8 5 12
rect 22 1 26 5
rect 44 1 48 5
rect 67 1 71 5
rect 96 1 100 5
rect 120 1 124 5
rect 149 1 153 5
rect 173 1 177 5
rect 202 1 206 5
rect 226 1 230 5
rect 256 1 260 5
rect 279 1 283 5
rect 309 1 313 5
rect 332 1 336 5
rect 361 1 365 5
rect 385 1 389 5
rect 415 1 419 5
rect 438 1 442 5
<< metal3 >>
rect 0 696 6 697
rect 0 692 1 696
rect 5 692 6 696
rect 0 691 6 692
rect 0 618 6 619
rect 0 614 1 618
rect 5 614 6 618
rect 0 613 6 614
rect 0 568 6 569
rect 0 564 1 568
rect 5 564 6 568
rect 0 563 6 564
rect 0 488 6 489
rect 0 484 1 488
rect 5 484 6 488
rect 0 483 6 484
rect 0 437 6 438
rect 0 433 1 437
rect 5 433 6 437
rect 0 432 6 433
rect 0 358 6 359
rect 0 354 1 358
rect 5 354 6 358
rect 0 353 6 354
rect 0 307 6 308
rect 0 303 1 307
rect 5 303 6 307
rect 0 302 6 303
rect 0 228 6 229
rect 0 224 1 228
rect 5 224 6 228
rect 0 223 6 224
rect 0 177 6 178
rect 0 173 1 177
rect 5 173 6 177
rect 0 172 6 173
rect 0 110 6 111
rect 0 106 1 110
rect 5 106 6 110
rect 0 105 6 106
rect 0 12 6 13
rect 0 8 1 12
rect 5 8 6 12
rect 0 7 6 8
rect 21 5 27 6
rect 21 1 22 5
rect 26 1 27 5
rect 21 0 27 1
rect 43 5 49 6
rect 43 1 44 5
rect 48 1 49 5
rect 43 0 49 1
rect 66 5 72 6
rect 66 1 67 5
rect 71 1 72 5
rect 66 0 72 1
rect 95 5 101 6
rect 95 1 96 5
rect 100 1 101 5
rect 95 0 101 1
rect 119 5 125 6
rect 119 1 120 5
rect 124 1 125 5
rect 119 0 125 1
rect 148 5 154 6
rect 148 1 149 5
rect 153 1 154 5
rect 148 0 154 1
rect 172 5 178 6
rect 172 1 173 5
rect 177 1 178 5
rect 172 0 178 1
rect 201 5 207 6
rect 201 1 202 5
rect 206 1 207 5
rect 201 0 207 1
rect 225 5 231 6
rect 225 1 226 5
rect 230 1 231 5
rect 225 0 231 1
rect 255 5 261 6
rect 255 1 256 5
rect 260 1 261 5
rect 255 0 261 1
rect 278 5 284 6
rect 278 1 279 5
rect 283 1 284 5
rect 278 0 284 1
rect 308 5 314 6
rect 308 1 309 5
rect 313 1 314 5
rect 308 0 314 1
rect 331 5 337 6
rect 331 1 332 5
rect 336 1 337 5
rect 331 0 337 1
rect 360 5 366 6
rect 360 1 361 5
rect 365 1 366 5
rect 360 0 366 1
rect 384 5 390 6
rect 384 1 385 5
rect 389 1 390 5
rect 384 0 390 1
rect 414 5 420 6
rect 414 1 415 5
rect 419 1 420 5
rect 414 0 420 1
rect 437 5 443 6
rect 437 1 438 5
rect 442 1 443 5
rect 437 0 443 1
<< labels >>
rlabel metal3 43 0 49 6 1 D[0]
rlabel metal3 66 0 72 6 1 Q[0]
rlabel metal3 95 0 101 6 1 D[1]
rlabel metal3 119 0 125 6 1 Q[1]
rlabel metal3 148 0 154 6 1 D[2]
rlabel metal3 172 0 178 6 1 Q[2]
rlabel metal3 201 0 207 6 1 D[3]
rlabel metal3 225 0 231 6 1 Q[3]
rlabel metal3 255 0 261 6 1 D[4]
rlabel metal3 278 0 284 6 1 Q[4]
rlabel metal3 308 0 314 6 1 D[5]
rlabel metal3 331 0 337 6 1 Q[5]
rlabel metal3 360 0 366 6 1 D[6]
rlabel metal3 384 0 390 6 1 Q[6]
rlabel metal3 414 0 420 6 1 D[7]
rlabel metal3 437 0 443 6 1 Q[7]
rlabel metal3 0 105 6 111 3 w
rlabel metal3 0 172 6 178 3 A[7]
rlabel metal3 0 223 6 229 3 A[6]
rlabel metal3 0 302 6 308 3 A[5]
rlabel metal3 0 353 6 359 3 A[4]
rlabel metal3 0 432 6 438 3 A[3]
rlabel metal3 0 483 6 489 3 A[2]
rlabel metal3 0 563 6 569 3 A[1]
rlabel metal3 0 613 6 619 3 A[0]
rlabel metal3 0 691 6 697 3 e
rlabel metal3 0 7 6 13 3 vdd
rlabel metal3 21 0 27 6 1 gnd
<< end >>

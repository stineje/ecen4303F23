# This is a template LEF file
# that can be used for a block macro
#
# Johannes Grad, IIT
#

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS


#########################################################
# CHANGE 1
# Change "SIZE" to the actual size of the block
# Currently the size is set to 138.9u wide, 213u high
#########################################################

SITE  MacroSite
    CLASS	Core ;
    SIZE	138.9 by 213 ;
END  MacroSite

#########################################################
# CHANGE 2
# Set SIZE to the same value as above
#########################################################

MACRO sram
  SIZE 138.9 by 213 ;
  CLASS BLOCK ;
  FOREIGN sram 0 0 ;
  ORIGIN 0 0 ;
  SYMMETRY x y r90 ;
  SITE MacroSite ;

#########################################################
# CHANGE 3
# Insert all the pin geometries
#########################################################

  Pin D[0]
    PORT
    LAYER metal3 ;
      RECT 12.9 0.0 14.7 1.8 ;
      END
  END D[0]

  Pin Q[0]
    PORT
    LAYER metal3 ;
      RECT 19.8 0.0 21.6 1.8 ;
      END
  END Q[0]

  Pin D[1]
    PORT
    LAYER metal3 ;
      RECT 28.5 0.0 30.3 1.8 ;
      END
  END D[1]

  Pin Q[1]
    PORT
    LAYER metal3 ;
      RECT 35.7 0.0 37.5 1.8 ;
      END
  END Q[1]

  Pin D[2]
    PORT
    LAYER metal3 ;
      RECT 44.4 0.0 46.2 1.8 ;
      END
  END D[2]

  Pin Q[2]
    PORT
    LAYER metal3 ;
      RECT 51.6 0.0 53.4 1.8 ;
      END
  END Q[2]

  Pin D[3]
    PORT
    LAYER metal3 ;
      RECT 60.3 0.0 62.1 1.8 ;
      END
  END D[3]

  Pin Q[3]
    PORT
    LAYER metal3 ;
      RECT 67.5 0.0 69.3 1.8 ;
      END
  END Q[3]

  Pin D[4]
    PORT
    LAYER metal3 ;
      RECT 76.5 0.0 78.3 1.8 ;
      END
  END D[4]

  Pin Q[4]
    PORT
    LAYER metal3 ;
      RECT 83.4 0.0 85.2 1.8 ;
      END
  END Q[4]

  Pin D[5]
    PORT
    LAYER metal3 ;
      RECT 92.4 0.0 94.2 1.8 ;
      END
  END D[5]

  Pin Q[5]
    PORT
    LAYER metal3 ;
      RECT 99.3 0.0 101.1 1.8 ;
      END
  END Q[5]

  Pin D[6]
    PORT
    LAYER metal3 ;
      RECT 108.0 0.0 109.8 1.8 ;
      END
  END D[6]

  Pin Q[6]
    PORT
    LAYER metal3 ;
      RECT 115.2 0.0 117.0 1.8 ;
      END
  END Q[6]

  Pin D[7]
    PORT
    LAYER metal3 ;
      RECT 124.2 0.0 126.0 1.8 ;
      END
  END D[7]

  Pin Q[7]
    PORT
    LAYER metal3 ;
      RECT 131.1 0.0 132.9 1.8 ;
      END
  END Q[7]

  Pin w
    PORT
    LAYER metal3 ;
      RECT 0.0 31.5 1.8 33.3 ;
      END
  END w

  Pin A[7]
    PORT
    LAYER metal3 ;
      RECT 0.0 51.6 1.8 53.4 ;
      END
  END A[7]

  Pin A[6]
    PORT
    LAYER metal3 ;
      RECT 0.0 66.9 1.8 68.7 ;
      END
  END A[6]

  Pin A[5]
    PORT
    LAYER metal3 ;
      RECT 0.0 90.6 1.8 92.4 ;
      END
  END A[5]

  Pin A[4]
    PORT
    LAYER metal3 ;
      RECT 0.0 105.9 1.8 107.7 ;
      END
  END A[4]

  Pin A[3]
    PORT
    LAYER metal3 ;
      RECT 0.0 129.6 1.8 131.4 ;
      END
  END A[3]

  Pin A[2]
    PORT
    LAYER metal3 ;
      RECT 0.0 144.9 1.8 146.7 ;
      END
  END A[2]

  Pin A[1]
    PORT
    LAYER metal3 ;
      RECT 0.0 168.9 1.8 170.7 ;
      END
  END A[1]

  Pin A[0]
    PORT
    LAYER metal3 ;
      RECT 0.0 183.9 1.8 185.7 ;
      END
  END A[0]

  Pin e
    PORT
    LAYER metal3 ;
      RECT 0.0 207.3 1.8 209.1 ;
      END
  END e

  Pin vdd
    USE POWER ;
    PORT
    LAYER metal3 ;
      RECT 0.0 2.1 1.8 3.9 ;
      END
  END vdd

  Pin gnd
    USE GROUND ;
    PORT
    LAYER metal3 ;
      RECT 6.3 0.0 8.1 1.8 ;
      END
  END gnd
 
#########################################################
# CHANGE 4
# Give lower left and upper right corner of obstruction
# metal1 and metal2 should cover the entire cell
# metal3 has to leave the pin area exposed
#########################################################

  OBS 
      LAYER metal1 ;
        RECT 0.0 0.0 138.9 213 ;
      LAYER metal2 ;
        RECT 0.0 0.0 138.9 213 ;
#      LAYER metal3 ;
#        RECT 2.7 2.7 138.9 213 ;
  END 

END sram

END LIBRARY

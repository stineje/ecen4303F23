magic
tech scmos
timestamp 1091055161
<< hvnwell >>
rect 17 634 433 996
rect -3 376 453 493
rect -3 14 17 376
rect 433 14 453 376
rect -3 -3 453 14
<< hvpwell >>
rect -3 999 453 1013
rect -3 631 14 999
rect 436 631 453 999
rect -3 517 453 631
rect 17 14 433 376
<< hvpsubstratepdiff >>
rect 0 1009 450 1010
rect 449 1005 450 1009
rect 0 1002 450 1005
rect 0 1000 11 1002
rect 9 628 11 1000
rect 439 1000 450 1002
rect 439 628 440 1000
rect 9 626 440 628
rect 449 626 450 1000
rect 0 620 450 626
rect 0 616 1 620
rect 0 610 450 616
rect 0 606 1 610
rect 0 600 450 606
rect 0 596 1 600
rect 0 590 450 596
rect 0 586 1 590
rect 0 580 450 586
rect 0 576 1 580
rect 0 570 450 576
rect 0 566 1 570
rect 0 560 450 566
rect 0 556 1 560
rect 0 550 450 556
rect 0 546 1 550
rect 0 540 450 546
rect 0 536 1 540
rect 0 530 450 536
rect 0 526 1 530
rect 0 520 450 526
rect 20 372 430 373
rect 20 363 21 372
rect 425 363 430 372
rect 20 361 430 363
rect 20 357 22 361
rect 426 357 430 361
rect 20 351 430 357
rect 20 347 22 351
rect 426 347 430 351
rect 20 341 430 347
rect 20 337 22 341
rect 426 337 430 341
rect 20 331 430 337
rect 20 327 22 331
rect 426 327 430 331
rect 20 321 430 327
rect 20 317 22 321
rect 426 317 430 321
rect 20 311 430 317
rect 20 307 22 311
rect 426 307 430 311
rect 20 301 430 307
rect 20 297 22 301
rect 426 297 430 301
rect 20 291 430 297
rect 20 287 22 291
rect 426 287 430 291
rect 20 281 430 287
rect 20 277 22 281
rect 426 277 430 281
rect 20 271 430 277
rect 20 267 22 271
rect 426 267 430 271
rect 20 261 430 267
rect 20 257 22 261
rect 426 257 430 261
rect 20 251 430 257
rect 20 247 22 251
rect 426 247 430 251
rect 20 241 430 247
rect 20 237 22 241
rect 426 237 430 241
rect 20 231 430 237
rect 20 227 22 231
rect 426 227 430 231
rect 20 221 430 227
rect 20 217 22 221
rect 426 217 430 221
rect 20 211 430 217
rect 20 207 22 211
rect 426 207 430 211
rect 20 201 430 207
rect 20 197 22 201
rect 426 197 430 201
rect 20 191 430 197
rect 20 187 22 191
rect 426 187 430 191
rect 20 181 430 187
rect 20 172 22 181
rect 426 172 430 181
rect 20 166 430 172
rect 20 162 22 166
rect 426 162 430 166
rect 20 156 430 162
rect 20 152 22 156
rect 426 152 430 156
rect 20 146 430 152
rect 20 142 22 146
rect 426 142 430 146
rect 20 136 430 142
rect 20 132 22 136
rect 426 132 430 136
rect 20 126 430 132
rect 20 122 22 126
rect 426 122 430 126
rect 20 116 430 122
rect 20 112 22 116
rect 426 112 430 116
rect 20 106 430 112
rect 20 102 22 106
rect 426 102 430 106
rect 20 96 430 102
rect 20 92 22 96
rect 426 92 430 96
rect 20 86 430 92
rect 20 82 22 86
rect 426 82 430 86
rect 20 76 430 82
rect 20 72 22 76
rect 426 72 430 76
rect 20 66 430 72
rect 20 62 22 66
rect 426 62 430 66
rect 20 56 430 62
rect 20 52 22 56
rect 426 52 430 56
rect 20 46 430 52
rect 20 42 22 46
rect 426 42 430 46
rect 20 36 430 42
rect 20 32 22 36
rect 426 32 430 36
rect 20 26 430 32
rect 20 22 22 26
rect 426 22 430 26
rect 20 17 430 22
<< hvnsubstratendiff >>
rect 20 991 430 993
rect 20 987 23 991
rect 427 987 430 991
rect 20 981 430 987
rect 20 977 23 981
rect 427 977 430 981
rect 20 971 430 977
rect 20 967 23 971
rect 427 967 430 971
rect 20 961 430 967
rect 20 957 23 961
rect 427 957 430 961
rect 20 951 430 957
rect 20 947 23 951
rect 427 947 430 951
rect 20 941 430 947
rect 20 937 23 941
rect 427 937 430 941
rect 20 931 430 937
rect 20 927 23 931
rect 427 927 430 931
rect 20 921 430 927
rect 20 917 23 921
rect 427 917 430 921
rect 20 911 430 917
rect 20 907 23 911
rect 427 907 430 911
rect 20 901 430 907
rect 20 897 23 901
rect 427 897 430 901
rect 20 891 430 897
rect 20 887 23 891
rect 427 887 430 891
rect 20 881 430 887
rect 20 877 23 881
rect 427 877 430 881
rect 20 871 430 877
rect 20 867 23 871
rect 427 867 430 871
rect 20 861 430 867
rect 20 857 23 861
rect 427 857 430 861
rect 20 851 430 857
rect 20 847 23 851
rect 427 847 430 851
rect 20 841 430 847
rect 20 837 23 841
rect 427 837 430 841
rect 20 831 430 837
rect 20 827 23 831
rect 427 827 430 831
rect 20 821 430 827
rect 20 817 23 821
rect 427 817 430 821
rect 20 811 430 817
rect 20 807 23 811
rect 427 807 430 811
rect 20 801 430 807
rect 20 797 23 801
rect 427 797 430 801
rect 20 791 430 797
rect 20 787 23 791
rect 427 787 430 791
rect 20 781 430 787
rect 20 777 23 781
rect 427 777 430 781
rect 20 771 430 777
rect 20 767 23 771
rect 427 767 430 771
rect 20 761 430 767
rect 20 757 23 761
rect 427 757 430 761
rect 20 751 430 757
rect 20 747 23 751
rect 427 747 430 751
rect 20 741 430 747
rect 20 737 23 741
rect 427 737 430 741
rect 20 731 430 737
rect 20 727 23 731
rect 427 727 430 731
rect 20 721 430 727
rect 20 717 23 721
rect 427 717 430 721
rect 20 711 430 717
rect 20 707 23 711
rect 427 707 430 711
rect 20 701 430 707
rect 20 697 23 701
rect 427 697 430 701
rect 20 691 430 697
rect 20 687 23 691
rect 427 687 430 691
rect 20 681 430 687
rect 20 677 23 681
rect 427 677 430 681
rect 20 671 430 677
rect 20 667 23 671
rect 427 667 430 671
rect 20 661 430 667
rect 20 657 23 661
rect 427 657 430 661
rect 20 647 430 657
rect 20 638 23 647
rect 427 638 430 647
rect 20 637 430 638
rect 0 484 450 490
rect 449 480 450 484
rect 0 474 450 480
rect 449 470 450 474
rect 0 464 450 470
rect 449 460 450 464
rect 0 454 450 460
rect 449 450 450 454
rect 0 444 450 450
rect 449 440 450 444
rect 0 434 450 440
rect 449 430 450 434
rect 0 424 450 430
rect 449 420 450 424
rect 0 414 450 420
rect 449 410 450 414
rect 0 404 450 410
rect 449 400 450 404
rect 0 394 450 400
rect 449 390 450 394
rect 0 384 450 390
rect 0 380 12 384
rect 131 380 134 384
rect 318 380 320 384
rect 434 380 450 384
rect 0 379 450 380
rect 0 0 2 379
rect 11 11 13 379
rect 436 11 439 379
rect 11 9 439 11
rect 11 0 15 9
rect 159 0 163 9
rect 287 0 291 9
rect 435 0 439 9
rect 448 0 450 379
<< hvpsubstratepcontact >>
rect 0 1005 449 1009
rect 0 626 9 1000
rect 440 626 449 1000
rect 1 616 450 620
rect 1 606 450 610
rect 1 596 450 600
rect 1 586 450 590
rect 1 576 450 580
rect 1 566 450 570
rect 1 556 450 560
rect 1 546 450 550
rect 1 536 450 540
rect 1 526 450 530
rect 21 363 425 372
rect 22 357 426 361
rect 22 347 426 351
rect 22 337 426 341
rect 22 327 426 331
rect 22 317 426 321
rect 22 307 426 311
rect 22 297 426 301
rect 22 287 426 291
rect 22 277 426 281
rect 22 267 426 271
rect 22 257 426 261
rect 22 247 426 251
rect 22 237 426 241
rect 22 227 426 231
rect 22 217 426 221
rect 22 207 426 211
rect 22 197 426 201
rect 22 187 426 191
rect 22 172 426 181
rect 22 162 426 166
rect 22 152 426 156
rect 22 142 426 146
rect 22 132 426 136
rect 22 122 426 126
rect 22 112 426 116
rect 22 102 426 106
rect 22 92 426 96
rect 22 82 426 86
rect 22 72 426 76
rect 22 62 426 66
rect 22 52 426 56
rect 22 42 426 46
rect 22 32 426 36
rect 22 22 426 26
<< hvnsubstratencontact >>
rect 23 987 427 991
rect 23 977 427 981
rect 23 967 427 971
rect 23 957 427 961
rect 23 947 427 951
rect 23 937 427 941
rect 23 927 427 931
rect 23 917 427 921
rect 23 907 427 911
rect 23 897 427 901
rect 23 887 427 891
rect 23 877 427 881
rect 23 867 427 871
rect 23 857 427 861
rect 23 847 427 851
rect 23 837 427 841
rect 23 827 427 831
rect 23 817 427 821
rect 23 807 427 811
rect 23 797 427 801
rect 23 787 427 791
rect 23 777 427 781
rect 23 767 427 771
rect 23 757 427 761
rect 23 747 427 751
rect 23 737 427 741
rect 23 727 427 731
rect 23 717 427 721
rect 23 707 427 711
rect 23 697 427 701
rect 23 687 427 691
rect 23 677 427 681
rect 23 667 427 671
rect 23 657 427 661
rect 23 638 427 647
rect 0 480 449 484
rect 0 470 449 474
rect 0 460 449 464
rect 0 450 449 454
rect 0 440 449 444
rect 0 430 449 434
rect 0 420 449 424
rect 0 410 449 414
rect 0 400 449 404
rect 0 390 449 394
rect 12 380 131 384
rect 134 380 318 384
rect 320 380 434 384
rect 2 0 11 379
rect 15 0 159 9
rect 163 0 287 9
rect 291 0 435 9
rect 439 0 448 379
<< metal1 >>
rect 0 1009 450 1010
rect 449 1005 450 1009
rect 0 1003 450 1005
rect 0 1000 10 1003
rect 9 627 10 1000
rect 440 1000 450 1003
rect 21 991 429 992
rect 21 987 23 991
rect 427 987 429 991
rect 21 986 429 987
rect 21 982 23 986
rect 427 982 429 986
rect 21 981 429 982
rect 21 977 23 981
rect 427 977 429 981
rect 21 976 429 977
rect 21 972 23 976
rect 427 972 429 976
rect 21 971 429 972
rect 21 967 23 971
rect 427 967 429 971
rect 21 966 429 967
rect 21 962 23 966
rect 427 962 429 966
rect 21 961 429 962
rect 21 957 23 961
rect 427 957 429 961
rect 21 956 429 957
rect 21 952 23 956
rect 427 952 429 956
rect 21 951 429 952
rect 21 947 23 951
rect 427 947 429 951
rect 21 946 429 947
rect 21 942 23 946
rect 427 942 429 946
rect 21 941 429 942
rect 21 937 23 941
rect 427 937 429 941
rect 21 936 429 937
rect 21 932 23 936
rect 427 932 429 936
rect 21 931 429 932
rect 21 927 23 931
rect 427 927 429 931
rect 21 926 429 927
rect 21 922 23 926
rect 427 922 429 926
rect 21 921 429 922
rect 21 917 23 921
rect 427 917 429 921
rect 21 916 429 917
rect 21 912 23 916
rect 427 912 429 916
rect 21 911 429 912
rect 21 907 23 911
rect 427 907 429 911
rect 21 906 429 907
rect 21 902 23 906
rect 427 902 429 906
rect 21 901 429 902
rect 21 897 23 901
rect 427 897 429 901
rect 21 896 429 897
rect 21 892 23 896
rect 427 892 429 896
rect 21 891 429 892
rect 21 887 23 891
rect 427 887 429 891
rect 21 886 429 887
rect 21 882 23 886
rect 427 882 429 886
rect 21 881 429 882
rect 21 877 23 881
rect 427 877 429 881
rect 21 876 429 877
rect 21 872 23 876
rect 427 872 429 876
rect 21 871 429 872
rect 21 867 23 871
rect 427 867 429 871
rect 21 866 429 867
rect 21 862 23 866
rect 427 862 429 866
rect 21 861 429 862
rect 21 857 23 861
rect 427 857 429 861
rect 21 856 429 857
rect 21 852 23 856
rect 427 852 429 856
rect 21 851 429 852
rect 21 847 23 851
rect 427 847 429 851
rect 21 846 429 847
rect 21 842 23 846
rect 427 842 429 846
rect 21 841 429 842
rect 21 837 23 841
rect 427 837 429 841
rect 21 836 429 837
rect 21 832 23 836
rect 427 832 429 836
rect 21 831 429 832
rect 21 827 23 831
rect 427 827 429 831
rect 21 826 429 827
rect 21 822 23 826
rect 427 822 429 826
rect 21 821 429 822
rect 21 817 23 821
rect 427 817 429 821
rect 21 816 429 817
rect 21 812 23 816
rect 427 812 429 816
rect 21 811 429 812
rect 21 807 23 811
rect 427 807 429 811
rect 21 806 429 807
rect 21 802 23 806
rect 427 802 429 806
rect 21 801 429 802
rect 21 797 23 801
rect 427 797 429 801
rect 21 796 429 797
rect 21 792 23 796
rect 427 792 429 796
rect 21 791 429 792
rect 21 787 23 791
rect 427 787 429 791
rect 21 786 429 787
rect 21 782 23 786
rect 427 782 429 786
rect 21 781 429 782
rect 21 777 23 781
rect 427 777 429 781
rect 21 776 429 777
rect 21 772 23 776
rect 427 772 429 776
rect 21 771 429 772
rect 21 767 23 771
rect 427 767 429 771
rect 21 766 429 767
rect 21 762 23 766
rect 427 762 429 766
rect 21 761 429 762
rect 21 757 23 761
rect 427 757 429 761
rect 21 756 429 757
rect 21 752 23 756
rect 427 752 429 756
rect 21 751 429 752
rect 21 747 23 751
rect 427 747 429 751
rect 21 746 429 747
rect 21 742 23 746
rect 427 742 429 746
rect 21 741 429 742
rect 21 737 23 741
rect 427 737 429 741
rect 21 736 429 737
rect 21 732 23 736
rect 427 732 429 736
rect 21 731 429 732
rect 21 727 23 731
rect 427 727 429 731
rect 21 726 429 727
rect 21 722 23 726
rect 427 722 429 726
rect 21 721 429 722
rect 21 717 23 721
rect 427 717 429 721
rect 21 716 429 717
rect 21 712 23 716
rect 427 712 429 716
rect 21 711 429 712
rect 21 707 23 711
rect 427 707 429 711
rect 21 706 429 707
rect 21 702 23 706
rect 427 702 429 706
rect 21 701 429 702
rect 21 697 23 701
rect 427 697 429 701
rect 21 696 429 697
rect 21 692 23 696
rect 427 692 429 696
rect 21 691 429 692
rect 21 687 23 691
rect 427 687 429 691
rect 21 686 429 687
rect 21 682 23 686
rect 427 682 429 686
rect 21 681 429 682
rect 21 677 23 681
rect 427 677 429 681
rect 21 676 429 677
rect 21 672 23 676
rect 427 672 429 676
rect 21 671 429 672
rect 21 667 23 671
rect 427 667 429 671
rect 21 666 429 667
rect 21 662 23 666
rect 427 662 429 666
rect 21 661 429 662
rect 21 657 23 661
rect 427 657 429 661
rect 21 656 429 657
rect 21 652 23 656
rect 427 652 429 656
rect 21 647 429 652
rect 21 638 23 647
rect 427 638 429 647
rect 9 626 440 627
rect 449 626 450 1000
rect 0 625 450 626
rect 0 621 1 625
rect 0 620 450 621
rect 0 616 1 620
rect 0 615 450 616
rect 0 611 1 615
rect 0 610 450 611
rect 0 606 1 610
rect 0 605 450 606
rect 0 601 1 605
rect 0 600 450 601
rect 0 596 1 600
rect 0 595 450 596
rect 0 591 1 595
rect 0 590 450 591
rect 0 586 1 590
rect 0 585 450 586
rect 0 581 1 585
rect 0 580 450 581
rect 0 576 1 580
rect 0 575 450 576
rect 0 571 1 575
rect 0 570 450 571
rect 0 566 1 570
rect 0 565 450 566
rect 0 561 1 565
rect 0 560 450 561
rect 0 556 1 560
rect 0 555 450 556
rect 0 551 1 555
rect 0 550 450 551
rect 0 546 1 550
rect 0 545 450 546
rect 0 541 1 545
rect 0 540 450 541
rect 0 536 1 540
rect 0 535 450 536
rect 0 531 1 535
rect 0 530 450 531
rect 0 526 1 530
rect 0 525 450 526
rect 0 521 1 525
rect 449 485 450 489
rect 0 484 450 485
rect 449 480 450 484
rect 0 479 450 480
rect 449 475 450 479
rect 0 474 450 475
rect 449 470 450 474
rect 0 469 450 470
rect 449 465 450 469
rect 0 464 450 465
rect 449 460 450 464
rect 0 459 450 460
rect 449 455 450 459
rect 0 454 450 455
rect 449 450 450 454
rect 0 449 450 450
rect 449 445 450 449
rect 0 444 450 445
rect 449 440 450 444
rect 0 439 450 440
rect 449 435 450 439
rect 0 434 450 435
rect 449 430 450 434
rect 0 429 450 430
rect 449 425 450 429
rect 0 424 450 425
rect 449 420 450 424
rect 0 419 450 420
rect 449 415 450 419
rect 0 414 450 415
rect 449 410 450 414
rect 0 409 450 410
rect 449 405 450 409
rect 0 404 450 405
rect 449 400 450 404
rect 0 399 450 400
rect 449 395 450 399
rect 0 394 450 395
rect 449 390 450 394
rect 0 389 450 390
rect 449 385 450 389
rect 0 384 450 385
rect 0 380 12 384
rect 131 380 134 384
rect 318 380 320 384
rect 434 380 450 384
rect 0 379 450 380
rect 0 0 2 379
rect 11 11 13 379
rect 425 363 429 372
rect 21 361 429 363
rect 21 357 22 361
rect 426 357 429 361
rect 21 356 429 357
rect 21 352 22 356
rect 426 352 429 356
rect 21 351 429 352
rect 21 347 22 351
rect 426 347 429 351
rect 21 346 429 347
rect 21 342 22 346
rect 426 342 429 346
rect 21 341 429 342
rect 21 337 22 341
rect 426 337 429 341
rect 21 336 429 337
rect 21 332 22 336
rect 426 332 429 336
rect 21 331 429 332
rect 21 327 22 331
rect 426 327 429 331
rect 21 326 429 327
rect 21 322 22 326
rect 426 322 429 326
rect 21 321 429 322
rect 21 317 22 321
rect 426 317 429 321
rect 21 316 429 317
rect 21 312 22 316
rect 426 312 429 316
rect 21 311 429 312
rect 21 307 22 311
rect 426 307 429 311
rect 21 306 429 307
rect 21 302 22 306
rect 426 302 429 306
rect 21 301 429 302
rect 21 297 22 301
rect 426 297 429 301
rect 21 296 429 297
rect 21 292 22 296
rect 426 292 429 296
rect 21 291 429 292
rect 21 287 22 291
rect 426 287 429 291
rect 21 286 429 287
rect 21 282 22 286
rect 426 282 429 286
rect 21 281 429 282
rect 21 277 22 281
rect 426 277 429 281
rect 21 276 429 277
rect 21 272 22 276
rect 426 272 429 276
rect 21 271 429 272
rect 21 267 22 271
rect 426 267 429 271
rect 21 266 429 267
rect 21 262 22 266
rect 426 262 429 266
rect 21 261 429 262
rect 21 257 22 261
rect 426 257 429 261
rect 21 256 429 257
rect 21 252 22 256
rect 426 252 429 256
rect 21 251 429 252
rect 21 247 22 251
rect 426 247 429 251
rect 21 246 429 247
rect 21 242 22 246
rect 426 242 429 246
rect 21 241 429 242
rect 21 237 22 241
rect 426 237 429 241
rect 21 236 429 237
rect 21 232 22 236
rect 426 232 429 236
rect 21 231 429 232
rect 21 227 22 231
rect 426 227 429 231
rect 21 226 429 227
rect 21 222 22 226
rect 426 222 429 226
rect 21 221 429 222
rect 21 217 22 221
rect 426 217 429 221
rect 21 216 429 217
rect 21 212 22 216
rect 426 212 429 216
rect 21 211 429 212
rect 21 207 22 211
rect 426 207 429 211
rect 21 206 429 207
rect 21 202 22 206
rect 426 202 429 206
rect 21 201 429 202
rect 21 197 22 201
rect 426 197 429 201
rect 21 196 429 197
rect 21 192 22 196
rect 426 192 429 196
rect 21 191 429 192
rect 21 187 22 191
rect 426 187 429 191
rect 21 186 429 187
rect 21 182 22 186
rect 426 182 429 186
rect 21 181 429 182
rect 21 172 22 181
rect 426 172 429 181
rect 21 171 429 172
rect 21 167 22 171
rect 426 167 429 171
rect 21 166 429 167
rect 21 162 22 166
rect 426 162 429 166
rect 21 161 429 162
rect 21 157 22 161
rect 426 157 429 161
rect 21 156 429 157
rect 21 152 22 156
rect 426 152 429 156
rect 21 151 429 152
rect 21 147 22 151
rect 426 147 429 151
rect 21 146 429 147
rect 21 142 22 146
rect 426 142 429 146
rect 21 141 429 142
rect 21 137 22 141
rect 426 137 429 141
rect 21 136 429 137
rect 21 132 22 136
rect 426 132 429 136
rect 21 131 429 132
rect 21 127 22 131
rect 426 127 429 131
rect 21 126 429 127
rect 21 122 22 126
rect 426 122 429 126
rect 21 121 429 122
rect 21 117 22 121
rect 426 117 429 121
rect 21 116 429 117
rect 21 112 22 116
rect 426 112 429 116
rect 21 111 429 112
rect 21 107 22 111
rect 426 107 429 111
rect 21 106 429 107
rect 21 102 22 106
rect 426 102 429 106
rect 21 101 429 102
rect 21 97 22 101
rect 426 97 429 101
rect 21 96 429 97
rect 21 92 22 96
rect 426 92 429 96
rect 21 91 429 92
rect 21 87 22 91
rect 426 87 429 91
rect 21 86 429 87
rect 21 82 22 86
rect 426 82 429 86
rect 21 81 429 82
rect 21 77 22 81
rect 426 77 429 81
rect 21 76 429 77
rect 21 72 22 76
rect 426 72 429 76
rect 21 71 429 72
rect 21 67 22 71
rect 426 67 429 71
rect 21 66 429 67
rect 21 62 22 66
rect 426 62 429 66
rect 21 61 429 62
rect 21 57 22 61
rect 426 57 429 61
rect 21 56 429 57
rect 21 52 22 56
rect 426 52 429 56
rect 21 51 429 52
rect 21 47 22 51
rect 426 47 429 51
rect 21 46 429 47
rect 21 42 22 46
rect 426 42 429 46
rect 21 41 429 42
rect 21 37 22 41
rect 426 37 429 41
rect 21 36 429 37
rect 21 32 22 36
rect 426 32 429 36
rect 21 31 429 32
rect 21 27 22 31
rect 426 27 429 31
rect 21 26 429 27
rect 21 22 22 26
rect 426 22 429 26
rect 21 18 429 22
rect 436 11 439 379
rect 11 9 439 11
rect 11 0 15 9
rect 159 0 163 9
rect 287 0 291 9
rect 435 0 439 9
rect 448 0 450 379
<< m2contact >>
rect 23 982 427 986
rect 23 972 427 976
rect 23 962 427 966
rect 23 952 427 956
rect 23 942 427 946
rect 23 932 427 936
rect 23 922 427 926
rect 23 912 427 916
rect 23 902 427 906
rect 23 892 427 896
rect 23 882 427 886
rect 23 872 427 876
rect 23 862 427 866
rect 23 852 427 856
rect 23 842 427 846
rect 23 832 427 836
rect 23 822 427 826
rect 23 812 427 816
rect 23 802 427 806
rect 23 792 427 796
rect 23 782 427 786
rect 23 772 427 776
rect 23 762 427 766
rect 23 752 427 756
rect 23 742 427 746
rect 23 732 427 736
rect 23 722 427 726
rect 23 712 427 716
rect 23 702 427 706
rect 23 692 427 696
rect 23 682 427 686
rect 23 672 427 676
rect 23 662 427 666
rect 23 652 427 656
rect 1 621 450 625
rect 1 611 450 615
rect 1 601 450 605
rect 1 591 450 595
rect 1 581 450 585
rect 1 571 450 575
rect 1 561 450 565
rect 1 551 450 555
rect 1 541 450 545
rect 1 531 450 535
rect 1 521 450 525
rect 0 485 449 489
rect 0 475 449 479
rect 0 465 449 469
rect 0 455 449 459
rect 0 445 449 449
rect 0 435 449 439
rect 0 425 449 429
rect 0 415 449 419
rect 0 405 449 409
rect 0 395 449 399
rect 0 385 449 389
rect 22 352 426 356
rect 22 342 426 346
rect 22 332 426 336
rect 22 322 426 326
rect 22 312 426 316
rect 22 302 426 306
rect 22 292 426 296
rect 22 282 426 286
rect 22 272 426 276
rect 22 262 426 266
rect 22 252 426 256
rect 22 242 426 246
rect 22 232 426 236
rect 22 222 426 226
rect 22 212 426 216
rect 22 202 426 206
rect 22 192 426 196
rect 22 182 426 186
rect 22 167 426 171
rect 22 157 426 161
rect 22 147 426 151
rect 22 137 426 141
rect 22 127 426 131
rect 22 117 426 121
rect 22 107 426 111
rect 22 97 426 101
rect 22 87 426 91
rect 22 77 426 81
rect 22 67 426 71
rect 22 57 426 61
rect 22 47 426 51
rect 22 37 426 41
rect 22 27 426 31
<< metal2 >>
rect 0 986 450 1010
rect 0 982 23 986
rect 427 982 450 986
rect 0 976 450 982
rect 0 972 23 976
rect 427 972 450 976
rect 0 966 450 972
rect 0 962 23 966
rect 427 962 450 966
rect 0 956 450 962
rect 0 952 23 956
rect 427 952 450 956
rect 0 946 450 952
rect 0 942 23 946
rect 427 942 450 946
rect 0 936 450 942
rect 0 932 23 936
rect 427 932 450 936
rect 0 926 450 932
rect 0 922 23 926
rect 427 922 450 926
rect 0 916 450 922
rect 0 912 23 916
rect 427 912 450 916
rect 0 906 450 912
rect 0 902 23 906
rect 427 902 450 906
rect 0 896 450 902
rect 0 892 23 896
rect 427 892 450 896
rect 0 886 450 892
rect 0 882 23 886
rect 427 882 450 886
rect 0 876 450 882
rect 0 872 23 876
rect 427 872 450 876
rect 0 866 450 872
rect 0 862 23 866
rect 427 862 450 866
rect 0 856 450 862
rect 0 852 23 856
rect 427 852 450 856
rect 0 846 450 852
rect 0 842 23 846
rect 427 842 450 846
rect 0 836 450 842
rect 0 832 23 836
rect 427 832 450 836
rect 0 826 450 832
rect 0 822 23 826
rect 427 822 450 826
rect 0 816 450 822
rect 0 812 23 816
rect 427 812 450 816
rect 0 806 450 812
rect 0 802 23 806
rect 427 802 450 806
rect 0 796 450 802
rect 0 792 23 796
rect 427 792 450 796
rect 0 786 450 792
rect 0 782 23 786
rect 427 782 450 786
rect 0 776 450 782
rect 0 772 23 776
rect 427 772 450 776
rect 0 766 450 772
rect 0 762 23 766
rect 427 762 450 766
rect 0 756 450 762
rect 0 752 23 756
rect 427 752 450 756
rect 0 746 450 752
rect 0 742 23 746
rect 427 742 450 746
rect 0 736 450 742
rect 0 732 23 736
rect 427 732 450 736
rect 0 726 450 732
rect 0 722 23 726
rect 427 722 450 726
rect 0 716 450 722
rect 0 712 23 716
rect 427 712 450 716
rect 0 706 450 712
rect 0 702 23 706
rect 427 702 450 706
rect 0 696 450 702
rect 0 692 23 696
rect 427 692 450 696
rect 0 686 450 692
rect 0 682 23 686
rect 427 682 450 686
rect 0 676 450 682
rect 0 672 23 676
rect 427 672 450 676
rect 0 666 450 672
rect 0 662 23 666
rect 427 662 450 666
rect 0 656 450 662
rect 0 652 23 656
rect 427 652 450 656
rect 0 648 450 652
rect 0 625 450 626
rect 0 621 1 625
rect 0 615 450 621
rect 0 611 1 615
rect 0 605 450 611
rect 0 601 1 605
rect 0 595 450 601
rect 0 591 1 595
rect 0 585 450 591
rect 0 581 1 585
rect 0 575 450 581
rect 0 571 1 575
rect 0 565 450 571
rect 0 561 1 565
rect 0 555 450 561
rect 0 551 1 555
rect 0 545 450 551
rect 0 541 1 545
rect 0 535 450 541
rect 0 531 1 535
rect 0 525 450 531
rect 0 521 1 525
rect 449 485 450 489
rect 0 479 450 485
rect 449 475 450 479
rect 0 469 450 475
rect 449 465 450 469
rect 0 459 450 465
rect 449 455 450 459
rect 0 449 450 455
rect 449 445 450 449
rect 0 439 450 445
rect 449 435 450 439
rect 0 429 450 435
rect 449 425 450 429
rect 0 419 450 425
rect 449 415 450 419
rect 0 409 450 415
rect 449 405 450 409
rect 0 399 450 405
rect 449 395 450 399
rect 0 389 450 395
rect 449 385 450 389
rect 0 384 450 385
rect 0 356 450 362
rect 0 352 22 356
rect 426 352 450 356
rect 0 346 450 352
rect 0 342 22 346
rect 426 342 450 346
rect 0 336 450 342
rect 0 332 22 336
rect 426 332 450 336
rect 0 326 450 332
rect 0 322 22 326
rect 426 322 450 326
rect 0 316 450 322
rect 0 312 22 316
rect 426 312 450 316
rect 0 306 450 312
rect 0 302 22 306
rect 426 302 450 306
rect 0 296 450 302
rect 0 292 22 296
rect 426 292 450 296
rect 0 286 450 292
rect 0 282 22 286
rect 426 282 450 286
rect 0 276 450 282
rect 0 272 22 276
rect 426 272 450 276
rect 0 266 450 272
rect 0 262 22 266
rect 426 262 450 266
rect 0 256 450 262
rect 0 252 22 256
rect 426 252 450 256
rect 0 246 450 252
rect 0 242 22 246
rect 426 242 450 246
rect 0 236 450 242
rect 0 232 22 236
rect 426 232 450 236
rect 0 226 450 232
rect 0 222 22 226
rect 426 222 450 226
rect 0 216 450 222
rect 0 212 22 216
rect 426 212 450 216
rect 0 206 450 212
rect 0 202 22 206
rect 426 202 450 206
rect 0 196 450 202
rect 0 192 22 196
rect 426 192 450 196
rect 0 186 450 192
rect 0 182 22 186
rect 426 182 450 186
rect 0 171 450 182
rect 0 167 22 171
rect 426 167 450 171
rect 0 161 450 167
rect 0 157 22 161
rect 426 157 450 161
rect 0 151 450 157
rect 0 147 22 151
rect 426 147 450 151
rect 0 141 450 147
rect 0 137 22 141
rect 426 137 450 141
rect 0 131 450 137
rect 0 127 22 131
rect 426 127 450 131
rect 0 121 450 127
rect 0 117 22 121
rect 426 117 450 121
rect 0 111 450 117
rect 0 107 22 111
rect 426 107 450 111
rect 0 101 450 107
rect 0 97 22 101
rect 426 97 450 101
rect 0 91 450 97
rect 0 87 22 91
rect 426 87 450 91
rect 0 81 450 87
rect 0 77 22 81
rect 426 77 450 81
rect 0 71 450 77
rect 0 67 22 71
rect 426 67 450 71
rect 0 61 450 67
rect 0 57 22 61
rect 426 57 450 61
rect 0 51 450 57
rect 0 47 22 51
rect 426 47 450 51
rect 0 41 450 47
rect 0 37 22 41
rect 426 37 450 41
rect 0 31 450 37
rect 0 27 22 31
rect 426 27 450 31
rect 0 0 450 27
<< end >>

magic
tech sky130A
timestamp 1605719121
<< nsubdiff >>
rect 0 17 17 29
rect 0 -12 17 0
<< nsubdiffcont >>
rect 0 0 17 17
<< locali >>
rect -8 0 0 17
rect 17 0 25 17
<< end >>

magic
tech scmos
timestamp 1091055094
<< nwell >>
rect 30 1110 420 1500
<< hvnwell >>
rect 17 634 433 996
rect -3 378 453 493
rect -3 11 11 378
rect 439 11 453 378
rect -3 -3 453 11
<< hvpwell >>
rect -3 999 453 1013
rect -3 631 14 999
rect 436 631 453 999
rect -3 517 453 631
rect 11 11 439 378
<< hvntransistor >>
rect 38 345 213 348
rect 237 345 412 348
rect 38 284 213 287
rect 237 284 412 287
rect 38 263 213 266
rect 237 263 412 266
rect 38 203 213 206
rect 38 182 213 185
rect 237 203 412 206
rect 237 182 412 185
rect 38 122 213 125
rect 237 122 412 125
rect 38 101 213 104
rect 237 101 412 104
rect 38 41 213 44
rect 237 41 412 44
<< hvndiffusion >>
rect 38 356 213 357
rect 38 352 41 356
rect 170 352 213 356
rect 38 348 213 352
rect 38 321 213 345
rect 38 317 56 321
rect 195 317 213 321
rect 38 315 213 317
rect 38 311 56 315
rect 195 311 213 315
rect 38 287 213 311
rect 237 356 412 357
rect 237 352 280 356
rect 409 352 412 356
rect 237 348 412 352
rect 38 280 213 284
rect 38 276 41 280
rect 180 276 213 280
rect 38 274 213 276
rect 38 270 41 274
rect 180 270 213 274
rect 38 266 213 270
rect 237 321 412 345
rect 237 317 255 321
rect 394 317 412 321
rect 237 315 412 317
rect 237 311 255 315
rect 394 311 412 315
rect 237 287 412 311
rect 237 280 412 284
rect 237 276 270 280
rect 409 276 412 280
rect 237 274 412 276
rect 237 270 270 274
rect 409 270 412 274
rect 237 266 412 270
rect 38 239 213 263
rect 38 230 56 239
rect 195 230 213 239
rect 38 206 213 230
rect 38 199 213 203
rect 38 195 41 199
rect 180 195 213 199
rect 38 193 213 195
rect 38 189 41 193
rect 180 189 213 193
rect 38 185 213 189
rect 38 158 213 182
rect 38 149 56 158
rect 195 149 213 158
rect 38 125 213 149
rect 237 239 412 263
rect 237 230 255 239
rect 394 230 412 239
rect 237 206 412 230
rect 237 199 412 203
rect 237 195 270 199
rect 409 195 412 199
rect 237 193 412 195
rect 237 189 270 193
rect 409 189 412 193
rect 237 185 412 189
rect 237 158 412 182
rect 237 149 255 158
rect 394 149 412 158
rect 237 125 412 149
rect 38 118 213 122
rect 38 114 41 118
rect 180 114 213 118
rect 38 112 213 114
rect 38 108 41 112
rect 180 108 213 112
rect 38 104 213 108
rect 38 77 213 101
rect 38 68 56 77
rect 195 68 213 77
rect 38 44 213 68
rect 237 118 412 122
rect 237 114 270 118
rect 409 114 412 118
rect 237 112 412 114
rect 237 108 270 112
rect 409 108 412 112
rect 237 104 412 108
rect 38 37 213 41
rect 38 33 41 37
rect 170 33 213 37
rect 38 32 213 33
rect 237 77 412 101
rect 237 68 255 77
rect 394 68 412 77
rect 237 44 412 68
rect 237 37 412 41
rect 237 33 280 37
rect 409 33 412 37
rect 237 32 412 33
<< hvndcontact >>
rect 41 352 170 356
rect 56 317 195 321
rect 56 311 195 315
rect 280 352 409 356
rect 41 276 180 280
rect 41 270 180 274
rect 255 317 394 321
rect 255 311 394 315
rect 270 276 409 280
rect 270 270 409 274
rect 56 230 195 239
rect 41 195 180 199
rect 41 189 180 193
rect 56 149 195 158
rect 255 230 394 239
rect 270 195 409 199
rect 270 189 409 193
rect 255 149 394 158
rect 41 114 180 118
rect 41 108 180 112
rect 56 68 195 77
rect 270 114 409 118
rect 270 108 409 112
rect 41 33 170 37
rect 255 68 394 77
rect 280 33 409 37
<< hvpsubstratepdiff >>
rect 0 626 1 1010
rect 10 1009 450 1010
rect 10 1005 15 1009
rect 174 1005 276 1009
rect 435 1007 450 1009
rect 435 1005 440 1007
rect 10 1002 440 1005
rect 10 628 11 1002
rect 439 628 440 1002
rect 449 628 450 1007
rect 10 626 450 628
rect 0 621 450 626
rect 0 620 218 621
rect 0 616 3 620
rect 132 616 218 620
rect 0 612 218 616
rect 232 620 450 621
rect 232 616 318 620
rect 447 616 450 620
rect 232 612 450 616
rect 0 610 450 612
rect 0 606 3 610
rect 132 606 318 610
rect 447 606 450 610
rect 0 602 218 606
rect 232 602 450 606
rect 0 600 450 602
rect 0 596 3 600
rect 132 596 318 600
rect 447 596 450 600
rect 0 592 218 596
rect 232 592 450 596
rect 0 590 450 592
rect 0 586 3 590
rect 132 586 318 590
rect 447 586 450 590
rect 0 580 218 586
rect 0 576 3 580
rect 132 576 218 580
rect 0 570 218 576
rect 0 566 3 570
rect 132 566 218 570
rect 0 560 218 566
rect 0 556 3 560
rect 132 556 218 560
rect 0 552 218 556
rect 232 580 450 586
rect 232 576 318 580
rect 447 576 450 580
rect 232 570 450 576
rect 232 566 318 570
rect 447 566 450 570
rect 232 560 450 566
rect 232 556 318 560
rect 447 556 450 560
rect 232 552 450 556
rect 0 550 450 552
rect 0 546 3 550
rect 132 546 318 550
rect 447 546 450 550
rect 0 542 218 546
rect 232 542 450 546
rect 0 540 450 542
rect 0 536 3 540
rect 132 536 318 540
rect 447 536 450 540
rect 0 532 218 536
rect 232 532 450 536
rect 0 530 450 532
rect 0 526 3 530
rect 132 526 318 530
rect 447 526 450 530
rect 0 522 218 526
rect 232 522 450 526
rect 0 520 450 522
rect 14 374 436 375
rect 173 373 436 374
rect 173 365 277 373
rect 14 364 277 365
rect 14 360 436 364
rect 14 31 20 360
rect 24 359 426 360
rect 24 31 30 359
rect 38 357 213 359
rect 218 342 232 359
rect 237 357 412 359
rect 218 338 223 342
rect 227 338 232 342
rect 218 332 232 338
rect 218 323 223 332
rect 227 323 232 332
rect 218 317 232 323
rect 218 313 223 317
rect 227 313 232 317
rect 218 269 232 313
rect 218 265 223 269
rect 227 265 232 269
rect 218 259 232 265
rect 218 250 223 259
rect 227 250 232 259
rect 218 244 232 250
rect 218 235 223 244
rect 227 235 232 244
rect 218 229 232 235
rect 218 220 223 229
rect 227 220 232 229
rect 218 214 232 220
rect 218 210 223 214
rect 227 210 232 214
rect 218 172 232 210
rect 218 168 223 172
rect 227 168 232 172
rect 218 162 232 168
rect 218 153 223 162
rect 227 153 232 162
rect 218 147 232 153
rect 218 138 223 147
rect 227 138 232 147
rect 218 132 232 138
rect 218 123 223 132
rect 227 123 232 132
rect 218 117 232 123
rect 218 113 223 117
rect 227 113 232 117
rect 218 76 232 113
rect 218 72 223 76
rect 227 72 232 76
rect 218 66 232 72
rect 218 57 223 66
rect 227 57 232 66
rect 218 51 232 57
rect 218 47 223 51
rect 227 47 232 51
rect 14 30 30 31
rect 38 30 213 32
rect 218 30 232 47
rect 237 30 412 32
rect 14 29 412 30
rect 420 31 426 359
rect 430 31 436 360
rect 420 29 436 31
rect 14 24 436 29
rect 14 20 15 24
rect 169 20 281 24
rect 435 20 436 24
rect 14 14 436 20
<< hvnsubstratendiff >>
rect 20 991 430 993
rect 20 987 21 991
rect 20 981 430 987
rect 20 977 21 981
rect 20 971 430 977
rect 20 967 21 971
rect 20 961 430 967
rect 20 957 21 961
rect 20 951 430 957
rect 20 947 21 951
rect 20 941 430 947
rect 20 937 21 941
rect 20 931 430 937
rect 20 927 21 931
rect 20 921 430 927
rect 20 917 21 921
rect 20 911 430 917
rect 20 907 21 911
rect 20 901 430 907
rect 20 897 21 901
rect 20 891 430 897
rect 20 887 21 891
rect 20 881 430 887
rect 20 877 21 881
rect 20 871 430 877
rect 20 867 21 871
rect 20 861 430 867
rect 20 857 21 861
rect 20 851 430 857
rect 20 847 21 851
rect 20 841 430 847
rect 20 837 21 841
rect 20 831 430 837
rect 20 827 21 831
rect 20 821 430 827
rect 20 817 21 821
rect 20 811 430 817
rect 20 807 21 811
rect 20 801 430 807
rect 20 797 21 801
rect 20 791 430 797
rect 20 787 21 791
rect 20 781 430 787
rect 20 777 21 781
rect 20 771 430 777
rect 20 767 21 771
rect 20 761 430 767
rect 20 757 21 761
rect 20 751 430 757
rect 20 747 21 751
rect 20 741 430 747
rect 20 737 21 741
rect 20 731 430 737
rect 20 727 21 731
rect 20 721 430 727
rect 20 717 21 721
rect 20 711 430 717
rect 20 707 21 711
rect 20 701 430 707
rect 20 697 21 701
rect 20 691 430 697
rect 20 687 21 691
rect 20 681 430 687
rect 20 677 21 681
rect 20 671 430 677
rect 20 667 21 671
rect 20 661 430 667
rect 20 657 21 661
rect 20 647 430 657
rect 20 638 23 647
rect 427 638 430 647
rect 20 637 430 638
rect 0 483 450 490
rect 0 479 3 483
rect 447 479 450 483
rect 0 473 450 479
rect 0 469 3 473
rect 447 469 450 473
rect 0 463 450 469
rect 0 459 3 463
rect 447 459 450 463
rect 0 453 450 459
rect 0 449 3 453
rect 447 449 450 453
rect 0 443 450 449
rect 0 439 3 443
rect 447 439 450 443
rect 0 433 450 439
rect 0 429 3 433
rect 447 429 450 433
rect 0 423 450 429
rect 0 419 3 423
rect 447 419 450 423
rect 0 413 450 419
rect 0 409 3 413
rect 447 409 450 413
rect 0 403 450 409
rect 0 399 3 403
rect 447 399 450 403
rect 0 393 450 399
rect 0 389 3 393
rect 447 389 450 393
rect 0 381 450 389
rect 0 2 2 381
rect 6 8 8 381
rect 442 8 444 381
rect 6 6 444 8
rect 6 2 10 6
rect 149 2 153 6
rect 297 2 301 6
rect 440 2 444 6
rect 448 2 450 381
rect 0 0 450 2
<< hvpsubstratepcontact >>
rect 1 626 10 1010
rect 15 1005 174 1009
rect 276 1005 435 1009
rect 440 628 449 1007
rect 3 616 132 620
rect 218 612 232 621
rect 318 616 447 620
rect 3 606 132 610
rect 318 606 447 610
rect 218 602 232 606
rect 3 596 132 600
rect 318 596 447 600
rect 218 592 232 596
rect 3 586 132 590
rect 318 586 447 590
rect 3 576 132 580
rect 3 566 132 570
rect 3 556 132 560
rect 218 552 232 586
rect 318 576 447 580
rect 318 566 447 570
rect 318 556 447 560
rect 3 546 132 550
rect 318 546 447 550
rect 218 542 232 546
rect 3 536 132 540
rect 318 536 447 540
rect 218 532 232 536
rect 3 526 132 530
rect 318 526 447 530
rect 218 522 232 526
rect 14 365 173 374
rect 277 364 436 373
rect 20 31 24 360
rect 223 338 227 342
rect 223 323 227 332
rect 223 313 227 317
rect 223 265 227 269
rect 223 250 227 259
rect 223 235 227 244
rect 223 220 227 229
rect 223 210 227 214
rect 223 168 227 172
rect 223 153 227 162
rect 223 138 227 147
rect 223 123 227 132
rect 223 113 227 117
rect 223 72 227 76
rect 223 57 227 66
rect 223 47 227 51
rect 426 31 430 360
rect 15 20 169 24
rect 281 20 435 24
<< hvnsubstratencontact >>
rect 21 987 430 991
rect 21 977 430 981
rect 21 967 430 971
rect 21 957 430 961
rect 21 947 430 951
rect 21 937 430 941
rect 21 927 430 931
rect 21 917 430 921
rect 21 907 430 911
rect 21 897 430 901
rect 21 887 430 891
rect 21 877 430 881
rect 21 867 430 871
rect 21 857 430 861
rect 21 847 430 851
rect 21 837 430 841
rect 21 827 430 831
rect 21 817 430 821
rect 21 807 430 811
rect 21 797 430 801
rect 21 787 430 791
rect 21 777 430 781
rect 21 767 430 771
rect 21 757 430 761
rect 21 747 430 751
rect 21 737 430 741
rect 21 727 430 731
rect 21 717 430 721
rect 21 707 430 711
rect 21 697 430 701
rect 21 687 430 691
rect 21 677 430 681
rect 21 667 430 671
rect 21 657 430 661
rect 23 638 427 647
rect 3 479 447 483
rect 3 469 447 473
rect 3 459 447 463
rect 3 449 447 453
rect 3 439 447 443
rect 3 429 447 433
rect 3 419 447 423
rect 3 409 447 413
rect 3 399 447 403
rect 3 389 447 393
rect 2 2 6 381
rect 10 2 149 6
rect 153 2 297 6
rect 301 2 440 6
rect 444 2 448 381
<< polysilicon >>
rect 31 346 38 348
rect 31 42 32 346
rect 36 345 38 346
rect 213 345 216 348
rect 36 287 37 345
rect 234 345 237 348
rect 412 346 419 348
rect 412 345 414 346
rect 36 284 38 287
rect 213 284 216 287
rect 36 266 37 284
rect 413 287 414 345
rect 234 284 237 287
rect 412 284 414 287
rect 36 263 38 266
rect 213 263 216 266
rect 413 266 414 284
rect 36 206 37 263
rect 234 263 237 266
rect 412 263 414 266
rect 36 203 38 206
rect 213 203 216 206
rect 36 185 37 203
rect 36 182 38 185
rect 213 182 216 185
rect 36 125 37 182
rect 413 206 414 263
rect 234 203 237 206
rect 412 203 414 206
rect 413 185 414 203
rect 234 182 237 185
rect 412 182 414 185
rect 36 122 38 125
rect 213 122 216 125
rect 413 125 414 182
rect 36 104 37 122
rect 234 122 237 125
rect 412 122 414 125
rect 36 101 38 104
rect 213 101 216 104
rect 36 44 37 101
rect 413 104 414 122
rect 234 101 237 104
rect 412 101 414 104
rect 36 42 38 44
rect 31 41 38 42
rect 213 41 216 44
rect 413 44 414 101
rect 234 41 237 44
rect 412 42 414 44
rect 418 42 419 346
rect 412 41 419 42
<< polycontact >>
rect 32 42 36 346
rect 414 42 418 346
<< metal1 >>
rect 30 1495 420 1500
rect 30 1114 34 1495
rect 415 1114 420 1495
rect 30 1110 420 1114
rect 137 1100 313 1110
rect 147 1090 303 1100
rect 157 1080 293 1090
rect 167 1070 283 1080
rect 0 626 1 1010
rect 10 1009 175 1010
rect 10 1005 15 1009
rect 174 1005 175 1009
rect 10 1003 175 1005
rect 178 998 272 1070
rect 275 1009 450 1010
rect 275 1005 276 1009
rect 435 1007 450 1009
rect 435 1005 440 1007
rect 275 1003 440 1005
rect 181 992 269 998
rect 21 991 430 992
rect 21 986 430 987
rect 21 981 430 982
rect 21 976 430 977
rect 21 971 430 972
rect 21 966 430 967
rect 21 961 430 962
rect 21 956 430 957
rect 21 951 430 952
rect 21 946 430 947
rect 21 941 430 942
rect 21 936 430 937
rect 21 931 430 932
rect 21 926 430 927
rect 21 921 430 922
rect 21 916 430 917
rect 21 911 430 912
rect 21 906 430 907
rect 21 901 430 902
rect 21 896 430 897
rect 21 891 430 892
rect 21 886 430 887
rect 21 881 430 882
rect 21 876 430 877
rect 21 871 430 872
rect 21 866 430 867
rect 21 861 430 862
rect 21 856 430 857
rect 21 851 430 852
rect 21 846 430 847
rect 21 841 430 842
rect 21 836 430 837
rect 21 831 430 832
rect 21 826 430 827
rect 21 821 430 822
rect 21 816 430 817
rect 21 811 430 812
rect 21 806 430 807
rect 21 801 430 802
rect 21 796 430 797
rect 21 791 430 792
rect 21 786 430 787
rect 21 781 430 782
rect 21 776 430 777
rect 21 771 430 772
rect 21 766 430 767
rect 21 761 430 762
rect 21 756 430 757
rect 21 751 430 752
rect 21 746 430 747
rect 21 741 430 742
rect 21 736 430 737
rect 21 731 430 732
rect 21 726 430 727
rect 21 721 430 722
rect 21 716 430 717
rect 21 711 430 712
rect 21 706 430 707
rect 21 701 430 702
rect 21 696 430 697
rect 21 691 430 692
rect 21 686 430 687
rect 21 681 430 682
rect 21 676 430 677
rect 21 671 430 672
rect 21 666 430 667
rect 21 661 430 662
rect 21 656 430 657
rect 21 647 429 652
rect 21 638 23 647
rect 427 638 429 647
rect 138 627 311 638
rect 449 628 450 1007
rect 440 627 450 628
rect 10 626 135 627
rect 0 625 135 626
rect 0 621 3 625
rect 132 621 135 625
rect 0 620 135 621
rect 0 616 3 620
rect 132 616 135 620
rect 0 615 135 616
rect 0 611 3 615
rect 132 611 135 615
rect 0 610 135 611
rect 0 606 3 610
rect 132 606 135 610
rect 0 605 135 606
rect 0 601 3 605
rect 132 601 135 605
rect 0 600 135 601
rect 0 596 3 600
rect 132 596 135 600
rect 0 595 135 596
rect 0 591 3 595
rect 132 591 135 595
rect 0 590 135 591
rect 0 586 3 590
rect 132 586 135 590
rect 0 585 135 586
rect 0 581 3 585
rect 132 581 135 585
rect 0 580 135 581
rect 0 576 3 580
rect 132 576 135 580
rect 0 575 135 576
rect 0 571 3 575
rect 132 571 135 575
rect 0 570 135 571
rect 0 566 3 570
rect 132 566 135 570
rect 0 565 135 566
rect 0 561 3 565
rect 132 561 135 565
rect 0 560 135 561
rect 0 556 3 560
rect 132 556 135 560
rect 0 555 135 556
rect 0 551 3 555
rect 132 551 135 555
rect 0 550 135 551
rect 0 546 3 550
rect 132 546 135 550
rect 0 545 135 546
rect 0 541 3 545
rect 132 541 135 545
rect 0 540 135 541
rect 0 536 3 540
rect 132 536 135 540
rect 0 535 135 536
rect 0 531 3 535
rect 132 531 135 535
rect 0 530 135 531
rect 0 526 3 530
rect 132 526 135 530
rect 0 525 135 526
rect 0 521 3 525
rect 132 521 135 525
rect 138 489 175 627
rect 178 489 215 627
rect 218 621 232 624
rect 218 611 232 612
rect 218 606 232 607
rect 218 601 232 602
rect 218 596 232 597
rect 218 591 232 592
rect 218 586 232 587
rect 218 551 232 552
rect 218 546 232 547
rect 218 541 232 542
rect 218 536 232 537
rect 218 531 232 532
rect 218 526 232 527
rect 218 521 232 522
rect 236 489 272 627
rect 275 489 311 627
rect 314 625 450 627
rect 314 621 318 625
rect 447 621 450 625
rect 314 620 450 621
rect 314 616 318 620
rect 447 616 450 620
rect 314 615 450 616
rect 314 611 318 615
rect 447 611 450 615
rect 314 610 450 611
rect 314 606 318 610
rect 447 606 450 610
rect 314 605 450 606
rect 314 601 318 605
rect 447 601 450 605
rect 314 600 450 601
rect 314 596 318 600
rect 447 596 450 600
rect 314 595 450 596
rect 314 591 318 595
rect 447 591 450 595
rect 314 590 450 591
rect 314 586 318 590
rect 447 586 450 590
rect 314 585 450 586
rect 314 581 318 585
rect 447 581 450 585
rect 314 580 450 581
rect 314 576 318 580
rect 447 576 450 580
rect 314 575 450 576
rect 314 571 318 575
rect 447 571 450 575
rect 314 570 450 571
rect 314 566 318 570
rect 447 566 450 570
rect 314 565 450 566
rect 314 561 318 565
rect 447 561 450 565
rect 314 560 450 561
rect 314 556 318 560
rect 447 556 450 560
rect 314 555 450 556
rect 314 551 318 555
rect 447 551 450 555
rect 314 550 450 551
rect 314 546 318 550
rect 447 546 450 550
rect 314 545 450 546
rect 314 541 318 545
rect 447 541 450 545
rect 314 540 450 541
rect 314 536 318 540
rect 447 536 450 540
rect 314 535 450 536
rect 314 531 318 535
rect 447 531 450 535
rect 314 530 450 531
rect 314 526 318 530
rect 447 526 450 530
rect 314 525 450 526
rect 314 521 318 525
rect 447 521 450 525
rect 0 488 450 489
rect 0 484 3 488
rect 447 484 450 488
rect 0 483 450 484
rect 0 479 3 483
rect 447 479 450 483
rect 0 478 450 479
rect 0 474 3 478
rect 447 474 450 478
rect 0 473 450 474
rect 0 469 3 473
rect 447 469 450 473
rect 0 468 450 469
rect 0 464 3 468
rect 447 464 450 468
rect 0 463 450 464
rect 0 459 3 463
rect 447 459 450 463
rect 0 458 450 459
rect 0 454 3 458
rect 447 454 450 458
rect 0 453 450 454
rect 0 449 3 453
rect 447 449 450 453
rect 0 448 450 449
rect 0 444 3 448
rect 447 444 450 448
rect 0 443 450 444
rect 0 439 3 443
rect 447 439 450 443
rect 0 438 450 439
rect 0 434 3 438
rect 447 434 450 438
rect 0 433 450 434
rect 0 429 3 433
rect 447 429 450 433
rect 0 428 450 429
rect 0 424 3 428
rect 447 424 450 428
rect 0 423 450 424
rect 0 419 3 423
rect 447 419 450 423
rect 0 418 450 419
rect 0 414 3 418
rect 447 414 450 418
rect 0 413 450 414
rect 0 409 3 413
rect 447 409 450 413
rect 0 408 450 409
rect 0 404 3 408
rect 447 404 450 408
rect 0 403 450 404
rect 0 399 3 403
rect 447 399 450 403
rect 0 398 450 399
rect 0 394 3 398
rect 447 394 450 398
rect 0 393 450 394
rect 0 389 3 393
rect 447 389 450 393
rect 0 388 450 389
rect 0 384 3 388
rect 447 384 450 388
rect 0 381 450 384
rect 0 2 2 381
rect 6 8 8 381
rect 14 374 174 375
rect 173 365 174 374
rect 14 360 174 365
rect 14 31 15 360
rect 19 31 20 360
rect 24 31 25 360
rect 29 356 174 360
rect 29 352 41 356
rect 170 352 174 356
rect 29 346 174 352
rect 29 42 32 346
rect 36 344 174 346
rect 36 320 39 344
rect 48 340 54 344
rect 173 340 174 344
rect 178 345 272 381
rect 178 337 220 345
rect 36 318 48 320
rect 36 314 39 318
rect 36 312 48 314
rect 36 288 39 312
rect 51 321 220 337
rect 51 317 56 321
rect 195 317 220 321
rect 51 315 220 317
rect 51 311 56 315
rect 195 311 220 315
rect 223 337 227 338
rect 223 332 227 333
rect 223 322 227 323
rect 223 317 227 318
rect 230 337 272 345
rect 276 373 436 375
rect 276 364 277 373
rect 276 360 436 364
rect 276 356 421 360
rect 276 352 280 356
rect 409 352 421 356
rect 276 346 421 352
rect 276 344 414 346
rect 276 340 277 344
rect 396 340 402 344
rect 230 321 399 337
rect 230 317 255 321
rect 394 317 399 321
rect 230 315 399 317
rect 51 310 220 311
rect 230 311 255 315
rect 394 311 399 315
rect 230 310 399 311
rect 51 295 399 310
rect 411 320 414 344
rect 402 318 414 320
rect 411 314 414 318
rect 402 312 414 314
rect 48 288 54 292
rect 178 288 185 292
rect 36 280 185 288
rect 36 276 41 280
rect 180 276 185 280
rect 36 274 185 276
rect 36 270 41 274
rect 180 270 185 274
rect 36 262 185 270
rect 36 238 39 262
rect 48 258 54 262
rect 178 258 185 262
rect 189 272 261 295
rect 189 255 220 272
rect 36 236 48 238
rect 36 207 39 236
rect 51 239 220 255
rect 51 230 56 239
rect 195 230 220 239
rect 51 214 220 230
rect 48 207 54 211
rect 178 207 185 211
rect 36 199 185 207
rect 36 195 41 199
rect 180 195 185 199
rect 36 193 185 195
rect 36 189 41 193
rect 180 189 185 193
rect 36 181 185 189
rect 36 157 39 181
rect 48 177 54 181
rect 178 177 185 181
rect 189 207 220 214
rect 223 264 227 265
rect 223 259 227 260
rect 223 249 227 250
rect 223 244 227 245
rect 223 234 227 235
rect 223 229 227 230
rect 223 219 227 220
rect 223 214 227 215
rect 230 255 261 272
rect 265 288 272 292
rect 396 288 402 292
rect 411 288 414 312
rect 265 280 414 288
rect 265 276 270 280
rect 409 276 414 280
rect 265 274 414 276
rect 265 270 270 274
rect 409 270 414 274
rect 265 262 414 270
rect 265 258 272 262
rect 396 258 402 262
rect 230 239 399 255
rect 230 230 255 239
rect 394 230 399 239
rect 230 214 399 230
rect 411 238 414 262
rect 402 236 414 238
rect 230 207 261 214
rect 189 175 261 207
rect 265 207 272 211
rect 396 207 402 211
rect 411 207 414 236
rect 265 199 414 207
rect 265 195 270 199
rect 409 195 414 199
rect 265 193 414 195
rect 265 189 270 193
rect 409 189 414 193
rect 265 181 414 189
rect 265 177 272 181
rect 396 177 402 181
rect 189 174 220 175
rect 36 155 48 157
rect 36 126 39 155
rect 51 158 220 174
rect 230 174 261 175
rect 51 149 56 158
rect 195 149 220 158
rect 51 133 220 149
rect 48 126 54 130
rect 178 126 185 130
rect 36 118 185 126
rect 36 114 41 118
rect 180 114 185 118
rect 36 112 185 114
rect 36 108 41 112
rect 180 108 185 112
rect 36 100 185 108
rect 36 71 39 100
rect 48 96 54 100
rect 178 96 185 100
rect 189 110 220 133
rect 223 167 227 168
rect 223 162 227 163
rect 223 152 227 153
rect 223 147 227 148
rect 223 137 227 138
rect 223 132 227 133
rect 223 122 227 123
rect 223 117 227 118
rect 230 158 399 174
rect 230 149 255 158
rect 394 149 399 158
rect 230 133 399 149
rect 411 157 414 181
rect 402 155 414 157
rect 230 110 261 133
rect 189 93 261 110
rect 265 126 272 130
rect 396 126 402 130
rect 411 126 414 155
rect 265 118 414 126
rect 265 114 270 118
rect 409 114 414 118
rect 265 112 414 114
rect 265 108 270 112
rect 409 108 414 112
rect 265 100 414 108
rect 265 96 272 100
rect 396 96 402 100
rect 36 69 48 71
rect 36 45 39 69
rect 51 79 399 93
rect 51 77 220 79
rect 51 68 56 77
rect 195 68 220 77
rect 230 77 399 79
rect 51 52 220 68
rect 48 45 54 49
rect 173 45 174 49
rect 36 42 174 45
rect 29 37 174 42
rect 29 33 41 37
rect 170 33 174 37
rect 29 31 174 33
rect 14 29 174 31
rect 14 25 15 29
rect 169 25 174 29
rect 14 24 174 25
rect 14 20 15 24
rect 169 20 174 24
rect 14 19 174 20
rect 14 15 15 19
rect 169 15 174 19
rect 14 14 174 15
rect 177 44 220 52
rect 223 71 227 72
rect 223 66 227 67
rect 223 56 227 57
rect 223 51 227 52
rect 230 68 255 77
rect 394 68 399 77
rect 230 52 399 68
rect 411 71 414 100
rect 402 69 414 71
rect 230 44 273 52
rect 177 29 273 44
rect 177 15 178 29
rect 272 15 273 29
rect 177 8 273 15
rect 276 45 277 49
rect 396 45 402 49
rect 411 45 414 69
rect 276 42 414 45
rect 418 42 421 346
rect 276 37 421 42
rect 276 33 280 37
rect 409 33 421 37
rect 276 31 421 33
rect 425 31 426 360
rect 430 31 431 360
rect 435 31 436 360
rect 276 29 436 31
rect 276 25 281 29
rect 435 25 436 29
rect 276 24 436 25
rect 276 20 281 24
rect 435 20 436 24
rect 276 19 436 20
rect 276 15 281 19
rect 435 15 436 19
rect 276 14 436 15
rect 442 8 444 381
rect 6 6 444 8
rect 6 2 10 6
rect 149 2 153 6
rect 297 2 301 6
rect 440 2 444 6
rect 448 2 450 381
rect 0 0 450 2
<< m2contact >>
rect 21 982 430 986
rect 21 972 430 976
rect 21 962 430 966
rect 21 952 430 956
rect 21 942 430 946
rect 21 932 430 936
rect 21 922 430 926
rect 21 912 430 916
rect 21 902 430 906
rect 21 892 430 896
rect 21 882 430 886
rect 21 872 430 876
rect 21 862 430 866
rect 21 852 430 856
rect 21 842 430 846
rect 21 832 430 836
rect 21 822 430 826
rect 21 812 430 816
rect 21 802 430 806
rect 21 792 430 796
rect 21 782 430 786
rect 21 772 430 776
rect 21 762 430 766
rect 21 752 430 756
rect 21 742 430 746
rect 21 732 430 736
rect 21 722 430 726
rect 21 712 430 716
rect 21 702 430 706
rect 21 692 430 696
rect 21 682 430 686
rect 21 672 430 676
rect 21 662 430 666
rect 21 652 430 656
rect 3 621 132 625
rect 3 611 132 615
rect 3 601 132 605
rect 3 591 132 595
rect 3 581 132 585
rect 3 571 132 575
rect 3 561 132 565
rect 3 551 132 555
rect 3 541 132 545
rect 3 531 132 535
rect 3 521 132 525
rect 218 607 232 611
rect 218 597 232 601
rect 218 587 232 591
rect 218 547 232 551
rect 218 537 232 541
rect 218 527 232 531
rect 318 621 447 625
rect 318 611 447 615
rect 318 601 447 605
rect 318 591 447 595
rect 318 581 447 585
rect 318 571 447 575
rect 318 561 447 565
rect 318 551 447 555
rect 318 541 447 545
rect 318 531 447 535
rect 318 521 447 525
rect 3 484 447 488
rect 3 474 447 478
rect 3 464 447 468
rect 3 454 447 458
rect 3 444 447 448
rect 3 434 447 438
rect 3 424 447 428
rect 3 414 447 418
rect 3 404 447 408
rect 3 394 447 398
rect 3 384 447 388
rect 15 31 19 360
rect 25 31 29 360
rect 39 320 48 344
rect 54 340 173 344
rect 39 314 48 318
rect 39 288 48 312
rect 223 333 227 337
rect 223 318 227 322
rect 277 340 396 344
rect 402 320 411 344
rect 402 314 411 318
rect 54 288 178 292
rect 39 238 48 262
rect 54 258 178 262
rect 39 207 48 236
rect 54 207 178 211
rect 39 157 48 181
rect 54 177 178 181
rect 223 260 227 264
rect 223 245 227 249
rect 223 230 227 234
rect 223 215 227 219
rect 272 288 396 292
rect 402 288 411 312
rect 272 258 396 262
rect 402 238 411 262
rect 272 207 396 211
rect 402 207 411 236
rect 272 177 396 181
rect 39 126 48 155
rect 54 126 178 130
rect 39 71 48 100
rect 54 96 178 100
rect 223 163 227 167
rect 223 148 227 152
rect 223 133 227 137
rect 223 118 227 122
rect 402 157 411 181
rect 272 126 396 130
rect 402 126 411 155
rect 272 96 396 100
rect 39 45 48 69
rect 54 45 173 49
rect 15 25 169 29
rect 15 15 169 19
rect 223 67 227 71
rect 223 52 227 56
rect 402 71 411 100
rect 178 15 272 29
rect 277 45 396 49
rect 402 45 411 69
rect 421 31 425 360
rect 431 31 435 360
rect 281 25 435 29
rect 281 15 435 19
<< metal2 >>
rect 30 1495 420 1500
rect 30 1114 34 1495
rect 415 1114 420 1495
rect 30 1110 420 1114
rect 0 986 450 1010
rect 0 982 21 986
rect 430 982 450 986
rect 0 976 450 982
rect 0 972 21 976
rect 430 972 450 976
rect 0 966 450 972
rect 0 962 21 966
rect 430 962 450 966
rect 0 956 450 962
rect 0 952 21 956
rect 430 952 450 956
rect 0 946 450 952
rect 0 942 21 946
rect 430 942 450 946
rect 0 936 450 942
rect 0 932 21 936
rect 430 932 450 936
rect 0 926 450 932
rect 0 922 21 926
rect 430 922 450 926
rect 0 916 450 922
rect 0 912 21 916
rect 430 912 450 916
rect 0 906 450 912
rect 0 902 21 906
rect 430 902 450 906
rect 0 896 450 902
rect 0 892 21 896
rect 430 892 450 896
rect 0 886 450 892
rect 0 882 21 886
rect 430 882 450 886
rect 0 876 450 882
rect 0 872 21 876
rect 430 872 450 876
rect 0 866 450 872
rect 0 862 21 866
rect 430 862 450 866
rect 0 856 450 862
rect 0 852 21 856
rect 430 852 450 856
rect 0 846 450 852
rect 0 842 21 846
rect 430 842 450 846
rect 0 836 450 842
rect 0 832 21 836
rect 430 832 450 836
rect 0 826 450 832
rect 0 822 21 826
rect 430 822 450 826
rect 0 816 450 822
rect 0 812 21 816
rect 430 812 450 816
rect 0 806 450 812
rect 0 802 21 806
rect 430 802 450 806
rect 0 796 450 802
rect 0 792 21 796
rect 430 792 450 796
rect 0 786 450 792
rect 0 782 21 786
rect 430 782 450 786
rect 0 776 450 782
rect 0 772 21 776
rect 430 772 450 776
rect 0 766 450 772
rect 0 762 21 766
rect 430 762 450 766
rect 0 756 450 762
rect 0 752 21 756
rect 430 752 450 756
rect 0 746 450 752
rect 0 742 21 746
rect 430 742 450 746
rect 0 736 450 742
rect 0 732 21 736
rect 430 732 450 736
rect 0 726 450 732
rect 0 722 21 726
rect 430 722 450 726
rect 0 716 450 722
rect 0 712 21 716
rect 430 712 450 716
rect 0 706 450 712
rect 0 702 21 706
rect 430 702 450 706
rect 0 696 450 702
rect 0 692 21 696
rect 430 692 450 696
rect 0 686 450 692
rect 0 682 21 686
rect 430 682 450 686
rect 0 676 450 682
rect 0 672 21 676
rect 430 672 450 676
rect 0 666 450 672
rect 0 662 21 666
rect 430 662 450 666
rect 0 656 450 662
rect 0 652 21 656
rect 430 652 450 656
rect 0 648 450 652
rect 0 625 450 626
rect 0 621 3 625
rect 132 621 318 625
rect 447 621 450 625
rect 0 615 450 621
rect 0 611 3 615
rect 132 611 318 615
rect 447 611 450 615
rect 0 607 218 611
rect 232 607 450 611
rect 0 605 450 607
rect 0 601 3 605
rect 132 601 318 605
rect 447 601 450 605
rect 0 597 218 601
rect 232 597 450 601
rect 0 595 450 597
rect 0 591 3 595
rect 132 591 318 595
rect 447 591 450 595
rect 0 587 218 591
rect 232 587 450 591
rect 0 585 450 587
rect 0 581 3 585
rect 132 581 318 585
rect 447 581 450 585
rect 0 575 450 581
rect 0 571 3 575
rect 132 571 318 575
rect 447 571 450 575
rect 0 565 450 571
rect 0 561 3 565
rect 132 561 318 565
rect 447 561 450 565
rect 0 555 450 561
rect 0 551 3 555
rect 132 551 318 555
rect 447 551 450 555
rect 0 547 218 551
rect 232 547 450 551
rect 0 545 450 547
rect 0 541 3 545
rect 132 541 318 545
rect 447 541 450 545
rect 0 537 218 541
rect 232 537 450 541
rect 0 535 450 537
rect 0 531 3 535
rect 132 531 318 535
rect 447 531 450 535
rect 0 527 218 531
rect 232 527 450 531
rect 0 525 450 527
rect 0 521 3 525
rect 132 521 318 525
rect 447 521 450 525
rect 0 488 450 489
rect 0 484 3 488
rect 447 484 450 488
rect 0 478 450 484
rect 0 474 3 478
rect 447 474 450 478
rect 0 468 450 474
rect 0 464 3 468
rect 447 464 450 468
rect 0 458 450 464
rect 0 454 3 458
rect 447 454 450 458
rect 0 448 450 454
rect 0 444 3 448
rect 447 444 450 448
rect 0 438 450 444
rect 0 434 3 438
rect 447 434 450 438
rect 0 428 450 434
rect 0 424 3 428
rect 447 424 450 428
rect 0 418 450 424
rect 0 414 3 418
rect 447 414 450 418
rect 0 408 450 414
rect 0 404 3 408
rect 447 404 450 408
rect 0 398 450 404
rect 0 394 3 398
rect 447 394 450 398
rect 0 388 450 394
rect 0 384 3 388
rect 447 384 450 388
rect 0 360 450 362
rect 0 31 15 360
rect 19 31 25 360
rect 29 344 421 360
rect 29 341 39 344
rect 29 337 32 341
rect 36 337 39 341
rect 29 331 39 337
rect 29 327 32 331
rect 36 327 39 331
rect 29 321 39 327
rect 29 317 32 321
rect 36 320 39 321
rect 48 340 54 344
rect 173 340 277 344
rect 396 340 402 344
rect 48 337 402 340
rect 48 333 223 337
rect 227 333 402 337
rect 48 322 402 333
rect 48 320 223 322
rect 36 318 223 320
rect 227 320 402 322
rect 411 341 421 344
rect 411 337 414 341
rect 418 337 421 341
rect 411 331 421 337
rect 411 327 414 331
rect 418 327 421 331
rect 411 321 421 327
rect 411 320 414 321
rect 227 318 414 320
rect 36 317 39 318
rect 29 314 39 317
rect 48 314 402 318
rect 411 317 414 318
rect 418 317 421 321
rect 411 314 421 317
rect 29 312 421 314
rect 29 311 39 312
rect 29 307 32 311
rect 36 307 39 311
rect 29 301 39 307
rect 29 297 32 301
rect 36 297 39 301
rect 29 291 39 297
rect 29 287 32 291
rect 36 288 39 291
rect 48 292 402 312
rect 48 288 54 292
rect 178 288 272 292
rect 396 288 402 292
rect 411 311 421 312
rect 411 307 414 311
rect 418 307 421 311
rect 411 301 421 307
rect 411 297 414 301
rect 418 297 421 301
rect 411 291 421 297
rect 411 288 414 291
rect 36 287 414 288
rect 418 287 421 291
rect 29 281 421 287
rect 29 277 32 281
rect 36 277 414 281
rect 418 277 421 281
rect 29 271 421 277
rect 29 267 32 271
rect 36 267 414 271
rect 418 267 421 271
rect 29 264 421 267
rect 29 262 223 264
rect 29 261 39 262
rect 29 257 32 261
rect 36 257 39 261
rect 29 251 39 257
rect 29 247 32 251
rect 36 247 39 251
rect 29 241 39 247
rect 29 237 32 241
rect 36 238 39 241
rect 48 258 54 262
rect 178 260 223 262
rect 227 262 421 264
rect 227 260 272 262
rect 178 258 272 260
rect 396 258 402 262
rect 48 249 402 258
rect 48 245 223 249
rect 227 245 402 249
rect 48 238 402 245
rect 411 261 421 262
rect 411 257 414 261
rect 418 257 421 261
rect 411 251 421 257
rect 411 247 414 251
rect 418 247 421 251
rect 411 241 421 247
rect 411 238 414 241
rect 36 237 414 238
rect 418 237 421 241
rect 29 236 421 237
rect 29 231 39 236
rect 29 227 32 231
rect 36 227 39 231
rect 29 221 39 227
rect 29 217 32 221
rect 36 217 39 221
rect 29 211 39 217
rect 29 207 32 211
rect 36 207 39 211
rect 48 234 402 236
rect 48 230 223 234
rect 227 230 402 234
rect 48 219 402 230
rect 48 215 223 219
rect 227 215 402 219
rect 48 211 402 215
rect 48 207 54 211
rect 178 207 272 211
rect 396 207 402 211
rect 411 231 421 236
rect 411 227 414 231
rect 418 227 421 231
rect 411 221 421 227
rect 411 217 414 221
rect 418 217 421 221
rect 411 211 421 217
rect 411 207 414 211
rect 418 207 421 211
rect 29 201 421 207
rect 29 197 32 201
rect 36 197 414 201
rect 418 197 421 201
rect 29 191 421 197
rect 29 187 32 191
rect 36 187 414 191
rect 418 187 421 191
rect 29 181 421 187
rect 29 177 32 181
rect 36 177 39 181
rect 29 171 39 177
rect 29 167 32 171
rect 36 167 39 171
rect 29 161 39 167
rect 29 157 32 161
rect 36 157 39 161
rect 48 177 54 181
rect 178 177 272 181
rect 396 177 402 181
rect 48 167 402 177
rect 48 163 223 167
rect 227 163 402 167
rect 48 157 402 163
rect 411 177 414 181
rect 418 177 421 181
rect 411 171 421 177
rect 411 167 414 171
rect 418 167 421 171
rect 411 161 421 167
rect 411 157 414 161
rect 418 157 421 161
rect 29 155 421 157
rect 29 151 39 155
rect 29 147 32 151
rect 36 147 39 151
rect 29 141 39 147
rect 29 137 32 141
rect 36 137 39 141
rect 29 131 39 137
rect 29 127 32 131
rect 36 127 39 131
rect 29 126 39 127
rect 48 152 402 155
rect 48 148 223 152
rect 227 148 402 152
rect 48 137 402 148
rect 48 133 223 137
rect 227 133 402 137
rect 48 130 402 133
rect 48 126 54 130
rect 178 126 272 130
rect 396 126 402 130
rect 411 151 421 155
rect 411 147 414 151
rect 418 147 421 151
rect 411 141 421 147
rect 411 137 414 141
rect 418 137 421 141
rect 411 131 421 137
rect 411 127 414 131
rect 418 127 421 131
rect 411 126 421 127
rect 29 122 421 126
rect 29 121 223 122
rect 29 117 32 121
rect 36 118 223 121
rect 227 121 421 122
rect 227 118 414 121
rect 36 117 414 118
rect 418 117 421 121
rect 29 111 421 117
rect 29 107 32 111
rect 36 107 414 111
rect 418 107 421 111
rect 29 101 421 107
rect 29 97 32 101
rect 36 100 414 101
rect 36 97 39 100
rect 29 91 39 97
rect 29 87 32 91
rect 36 87 39 91
rect 29 81 39 87
rect 29 77 32 81
rect 36 77 39 81
rect 29 71 39 77
rect 48 96 54 100
rect 178 96 272 100
rect 396 96 402 100
rect 48 71 402 96
rect 411 97 414 100
rect 418 97 421 101
rect 411 91 421 97
rect 411 87 414 91
rect 418 87 421 91
rect 411 81 421 87
rect 411 77 414 81
rect 418 77 421 81
rect 411 71 421 77
rect 29 67 32 71
rect 36 69 223 71
rect 36 67 39 69
rect 29 61 39 67
rect 29 57 32 61
rect 36 57 39 61
rect 29 51 39 57
rect 29 47 32 51
rect 36 47 39 51
rect 29 45 39 47
rect 48 67 223 69
rect 227 69 414 71
rect 227 67 402 69
rect 48 56 402 67
rect 48 52 223 56
rect 227 52 402 56
rect 48 49 402 52
rect 48 45 54 49
rect 173 45 277 49
rect 396 45 402 49
rect 411 67 414 69
rect 418 67 421 71
rect 411 61 421 67
rect 411 57 414 61
rect 418 57 421 61
rect 411 51 421 57
rect 411 47 414 51
rect 418 47 421 51
rect 411 45 421 47
rect 29 34 421 45
rect 29 31 172 34
rect 0 29 172 31
rect 278 31 421 34
rect 425 31 431 360
rect 435 31 450 360
rect 278 29 450 31
rect 0 25 15 29
rect 169 25 172 29
rect 0 19 172 25
rect 0 15 15 19
rect 169 15 172 19
rect 0 0 172 15
rect 177 15 178 29
rect 272 15 273 29
rect 177 0 273 15
rect 278 25 281 29
rect 435 25 450 29
rect 278 19 450 25
rect 278 15 281 19
rect 435 15 450 19
rect 278 0 450 15
<< pad >>
rect 34 1114 415 1495
<< m1p >>
rect 177 0 273 4
<< m4p >>
rect 211 1330 222 1342
<< labels >>
rlabel metal1 225 0 225 0 8 vdd
rlabel m4p 216 1336 216 1336 1 YPAD
<< end >>

magic
tech sky130A
timestamp 1605718463
<< metal1 >>
rect 0 26 26 29
rect 0 -3 26 0
<< via1 >>
rect 0 0 26 26
<< metal2 >>
rect 0 26 26 29
rect 0 -3 26 0
<< end >>

magic
tech scmos
timestamp 1084294447
<< nwell >>
rect 20 740 280 1000
rect 17 429 283 653
rect -3 248 303 330
rect -3 11 11 248
rect 289 11 303 248
rect -3 -3 303 11
<< pwell >>
rect -3 656 303 673
rect -3 426 14 656
rect 286 426 303 656
rect -3 340 303 426
rect 11 11 289 248
<< ntransistor >>
rect 38 216 138 219
rect 162 216 262 219
rect 38 171 138 174
rect 38 150 138 153
rect 162 171 262 174
rect 162 150 262 153
rect 38 106 138 109
rect 38 85 138 88
rect 162 106 262 109
rect 162 85 262 88
rect 38 41 138 44
rect 162 41 262 44
<< ndiffusion >>
rect 38 227 138 228
rect 38 223 41 227
rect 95 223 138 227
rect 38 219 138 223
rect 162 227 262 228
rect 162 223 205 227
rect 259 223 262 227
rect 162 219 262 223
rect 38 200 138 216
rect 38 196 56 200
rect 120 196 138 200
rect 38 194 138 196
rect 38 190 56 194
rect 120 190 138 194
rect 38 174 138 190
rect 38 167 138 171
rect 38 163 41 167
rect 120 163 138 167
rect 38 161 138 163
rect 38 157 41 161
rect 120 157 138 161
rect 38 153 138 157
rect 38 134 138 150
rect 38 125 56 134
rect 120 125 138 134
rect 38 109 138 125
rect 162 200 262 216
rect 162 196 180 200
rect 244 196 262 200
rect 162 194 262 196
rect 162 190 180 194
rect 244 190 262 194
rect 162 174 262 190
rect 162 167 262 171
rect 162 163 180 167
rect 259 163 262 167
rect 162 161 262 163
rect 162 157 180 161
rect 259 157 262 161
rect 162 153 262 157
rect 38 102 138 106
rect 38 98 41 102
rect 120 98 138 102
rect 38 96 138 98
rect 38 92 41 96
rect 120 92 138 96
rect 38 88 138 92
rect 38 69 138 85
rect 38 60 56 69
rect 120 60 138 69
rect 38 44 138 60
rect 162 134 262 150
rect 162 125 180 134
rect 244 125 262 134
rect 162 109 262 125
rect 162 102 262 106
rect 162 98 180 102
rect 259 98 262 102
rect 162 96 262 98
rect 162 92 180 96
rect 259 92 262 96
rect 162 88 262 92
rect 162 69 262 85
rect 162 60 180 69
rect 244 60 262 69
rect 162 44 262 60
rect 38 37 138 41
rect 38 33 41 37
rect 95 33 138 37
rect 38 32 138 33
rect 162 37 262 41
rect 162 33 205 37
rect 259 33 262 37
rect 162 32 262 33
<< ndcontact >>
rect 41 223 95 227
rect 205 223 259 227
rect 56 196 120 200
rect 56 190 120 194
rect 41 163 120 167
rect 41 157 120 161
rect 56 125 120 134
rect 180 196 244 200
rect 180 190 244 194
rect 180 163 259 167
rect 180 157 259 161
rect 41 98 120 102
rect 41 92 120 96
rect 56 60 120 69
rect 180 125 244 134
rect 180 98 259 102
rect 180 92 259 96
rect 180 60 244 69
rect 41 33 95 37
rect 205 33 259 37
<< psubstratepdiff >>
rect 0 669 300 670
rect 0 660 1 669
rect 95 660 204 669
rect 298 660 300 669
rect 0 659 300 660
rect 0 658 11 659
rect 0 424 1 658
rect 10 424 11 658
rect 289 658 300 659
rect 0 423 11 424
rect 289 424 290 658
rect 299 424 300 658
rect 289 423 300 424
rect 0 418 300 423
rect 0 414 143 418
rect 157 414 204 418
rect 298 414 300 418
rect 0 413 300 414
rect 0 409 2 413
rect 96 409 300 413
rect 0 408 300 409
rect 0 404 143 408
rect 157 404 204 408
rect 298 404 300 408
rect 0 403 300 404
rect 0 399 2 403
rect 96 399 300 403
rect 0 398 300 399
rect 0 394 143 398
rect 157 394 204 398
rect 298 394 300 398
rect 0 393 300 394
rect 0 389 2 393
rect 96 389 300 393
rect 0 388 300 389
rect 0 384 143 388
rect 157 384 204 388
rect 298 384 300 388
rect 0 383 300 384
rect 0 379 2 383
rect 96 379 300 383
rect 0 378 300 379
rect 0 374 143 378
rect 157 374 204 378
rect 298 374 300 378
rect 0 373 300 374
rect 0 369 2 373
rect 96 369 300 373
rect 0 368 300 369
rect 0 364 143 368
rect 157 364 204 368
rect 298 364 300 368
rect 0 363 300 364
rect 0 359 2 363
rect 96 359 300 363
rect 0 358 300 359
rect 0 354 143 358
rect 157 354 204 358
rect 298 354 300 358
rect 0 348 300 354
rect 0 344 2 348
rect 96 344 143 348
rect 157 344 204 348
rect 298 344 300 348
rect 0 343 300 344
rect 14 244 286 245
rect 14 241 202 244
rect 14 237 19 241
rect 98 237 202 241
rect 14 235 202 237
rect 281 235 286 244
rect 14 233 286 235
rect 14 29 24 233
rect 28 230 39 233
rect 28 30 30 230
rect 38 229 39 230
rect 98 230 202 233
rect 98 229 138 230
rect 38 228 138 229
rect 142 223 158 230
rect 142 219 145 223
rect 154 219 158 223
rect 162 229 202 230
rect 261 230 277 233
rect 261 229 262 230
rect 162 228 262 229
rect 142 215 158 219
rect 142 211 145 215
rect 154 211 158 215
rect 142 207 158 211
rect 142 203 145 207
rect 154 203 158 207
rect 142 135 158 203
rect 142 131 145 135
rect 154 131 158 135
rect 142 127 158 131
rect 142 123 145 127
rect 154 123 158 127
rect 142 63 158 123
rect 142 59 145 63
rect 154 59 158 63
rect 142 55 158 59
rect 142 51 145 55
rect 154 51 158 55
rect 142 47 158 51
rect 142 43 145 47
rect 154 43 158 47
rect 38 30 138 32
rect 142 39 158 43
rect 142 35 145 39
rect 154 35 158 39
rect 142 30 158 35
rect 162 30 262 32
rect 270 30 277 230
rect 28 29 277 30
rect 281 29 286 233
rect 14 27 286 29
rect 14 23 19 27
rect 98 23 202 27
rect 281 23 286 27
rect 14 14 286 23
<< nsubstratendiff >>
rect 20 649 280 650
rect 20 645 23 649
rect 277 645 280 649
rect 20 639 280 645
rect 20 635 23 639
rect 277 635 280 639
rect 20 629 280 635
rect 20 625 23 629
rect 277 625 280 629
rect 20 619 280 625
rect 20 615 23 619
rect 277 615 280 619
rect 20 609 280 615
rect 20 605 23 609
rect 277 605 280 609
rect 20 599 280 605
rect 20 595 23 599
rect 277 595 280 599
rect 20 589 280 595
rect 20 585 23 589
rect 277 585 280 589
rect 20 579 280 585
rect 20 575 23 579
rect 277 575 280 579
rect 20 569 280 575
rect 20 565 23 569
rect 277 565 280 569
rect 20 559 280 565
rect 20 555 23 559
rect 277 555 280 559
rect 20 549 280 555
rect 20 545 23 549
rect 277 545 280 549
rect 20 539 280 545
rect 20 535 23 539
rect 277 535 280 539
rect 20 529 280 535
rect 20 525 23 529
rect 277 525 280 529
rect 20 519 280 525
rect 20 515 23 519
rect 277 515 280 519
rect 20 509 280 515
rect 20 505 23 509
rect 277 505 280 509
rect 20 499 280 505
rect 20 495 23 499
rect 277 495 280 499
rect 20 489 280 495
rect 20 485 23 489
rect 277 485 280 489
rect 20 479 280 485
rect 20 475 23 479
rect 277 475 280 479
rect 20 469 280 475
rect 20 465 23 469
rect 277 465 280 469
rect 20 459 280 465
rect 20 455 23 459
rect 277 455 280 459
rect 20 449 280 455
rect 20 445 23 449
rect 277 445 280 449
rect 20 439 280 445
rect 20 435 23 439
rect 277 435 280 439
rect 20 432 280 435
rect 0 326 300 327
rect 0 322 3 326
rect 297 322 300 326
rect 0 316 300 322
rect 0 312 3 316
rect 297 312 300 316
rect 0 306 300 312
rect 0 302 3 306
rect 297 302 300 306
rect 0 296 300 302
rect 0 292 3 296
rect 297 292 300 296
rect 0 286 300 292
rect 0 282 3 286
rect 297 282 300 286
rect 0 276 300 282
rect 0 272 3 276
rect 297 272 300 276
rect 0 266 300 272
rect 0 262 3 266
rect 297 262 300 266
rect 0 256 300 262
rect 0 3 2 256
rect 6 8 8 256
rect 292 8 294 256
rect 6 7 294 8
rect 6 3 8 7
rect 92 3 203 7
rect 292 3 294 7
rect 298 3 300 256
rect 0 0 300 3
<< psubstratepcontact >>
rect 1 660 95 669
rect 204 660 298 669
rect 1 424 10 658
rect 290 424 299 658
rect 143 414 157 418
rect 204 414 298 418
rect 2 409 96 413
rect 143 404 157 408
rect 204 404 298 408
rect 2 399 96 403
rect 143 394 157 398
rect 204 394 298 398
rect 2 389 96 393
rect 143 384 157 388
rect 204 384 298 388
rect 2 379 96 383
rect 143 374 157 378
rect 204 374 298 378
rect 2 369 96 373
rect 143 364 157 368
rect 204 364 298 368
rect 2 359 96 363
rect 143 354 157 358
rect 204 354 298 358
rect 2 344 96 348
rect 143 344 157 348
rect 204 344 298 348
rect 19 237 98 241
rect 202 235 281 244
rect 24 29 28 233
rect 39 229 98 233
rect 145 219 154 223
rect 202 229 261 233
rect 145 211 154 215
rect 145 203 154 207
rect 145 131 154 135
rect 145 123 154 127
rect 145 59 154 63
rect 145 51 154 55
rect 145 43 154 47
rect 145 35 154 39
rect 277 29 281 233
rect 19 23 98 27
rect 202 23 281 27
<< nsubstratencontact >>
rect 23 645 277 649
rect 23 635 277 639
rect 23 625 277 629
rect 23 615 277 619
rect 23 605 277 609
rect 23 595 277 599
rect 23 585 277 589
rect 23 575 277 579
rect 23 565 277 569
rect 23 555 277 559
rect 23 545 277 549
rect 23 535 277 539
rect 23 525 277 529
rect 23 515 277 519
rect 23 505 277 509
rect 23 495 277 499
rect 23 485 277 489
rect 23 475 277 479
rect 23 465 277 469
rect 23 455 277 459
rect 23 445 277 449
rect 23 435 277 439
rect 3 322 297 326
rect 3 312 297 316
rect 3 302 297 306
rect 3 292 297 296
rect 3 282 297 286
rect 3 272 297 276
rect 3 262 297 266
rect 2 3 6 256
rect 8 252 292 256
rect 8 3 92 7
rect 203 3 292 7
rect 294 3 298 256
<< polysilicon >>
rect 31 217 38 219
rect 31 43 32 217
rect 36 216 38 217
rect 138 216 140 219
rect 36 174 37 216
rect 160 216 162 219
rect 262 217 269 219
rect 262 216 264 217
rect 36 171 38 174
rect 138 171 140 174
rect 36 153 37 171
rect 36 150 38 153
rect 138 150 140 153
rect 36 109 37 150
rect 263 174 264 216
rect 160 171 162 174
rect 262 171 264 174
rect 263 153 264 171
rect 160 150 162 153
rect 262 150 264 153
rect 36 106 38 109
rect 138 106 140 109
rect 36 88 37 106
rect 36 85 38 88
rect 138 85 140 88
rect 36 44 37 85
rect 263 109 264 150
rect 160 106 162 109
rect 262 106 264 109
rect 263 88 264 106
rect 160 85 162 88
rect 262 85 264 88
rect 36 43 38 44
rect 31 41 38 43
rect 138 41 140 44
rect 263 44 264 85
rect 160 41 162 44
rect 262 43 264 44
rect 268 43 269 217
rect 262 41 269 43
<< polycontact >>
rect 32 43 36 217
rect 264 43 268 217
<< metal1 >>
rect 20 997 280 1000
rect 20 743 23 997
rect 277 743 280 997
rect 20 740 280 743
rect 62 730 238 740
rect 72 720 228 730
rect 82 710 218 720
rect 92 700 208 710
rect 0 669 99 670
rect 0 660 1 669
rect 95 660 99 669
rect 0 659 99 660
rect 0 658 10 659
rect 0 424 1 658
rect 102 650 198 700
rect 201 669 300 670
rect 201 660 204 669
rect 298 660 300 669
rect 201 659 300 660
rect 289 658 300 659
rect 50 649 280 650
rect 21 645 23 649
rect 277 645 280 649
rect 21 644 280 645
rect 21 640 23 644
rect 277 640 280 644
rect 21 639 280 640
rect 21 635 23 639
rect 277 635 280 639
rect 21 634 280 635
rect 21 630 23 634
rect 277 630 280 634
rect 21 629 280 630
rect 21 625 23 629
rect 277 625 280 629
rect 21 624 280 625
rect 21 620 23 624
rect 277 620 280 624
rect 21 619 280 620
rect 21 615 23 619
rect 277 615 280 619
rect 21 614 280 615
rect 21 610 23 614
rect 277 610 280 614
rect 21 609 280 610
rect 21 605 23 609
rect 277 605 280 609
rect 21 604 280 605
rect 21 600 23 604
rect 277 600 280 604
rect 21 599 280 600
rect 21 595 23 599
rect 277 595 280 599
rect 21 594 280 595
rect 21 590 23 594
rect 277 590 280 594
rect 21 589 280 590
rect 21 585 23 589
rect 277 585 280 589
rect 21 584 280 585
rect 21 580 23 584
rect 277 580 280 584
rect 21 579 280 580
rect 21 575 23 579
rect 277 575 280 579
rect 21 574 280 575
rect 21 570 23 574
rect 277 570 280 574
rect 21 569 280 570
rect 21 565 23 569
rect 277 565 280 569
rect 21 564 280 565
rect 21 560 23 564
rect 277 560 280 564
rect 21 559 280 560
rect 21 555 23 559
rect 277 555 280 559
rect 21 554 280 555
rect 21 550 23 554
rect 277 550 280 554
rect 21 549 280 550
rect 21 545 23 549
rect 277 545 280 549
rect 21 544 280 545
rect 21 540 23 544
rect 277 540 280 544
rect 21 539 280 540
rect 21 535 23 539
rect 277 535 280 539
rect 21 534 280 535
rect 21 530 23 534
rect 277 530 280 534
rect 21 529 280 530
rect 21 525 23 529
rect 277 525 280 529
rect 21 524 280 525
rect 21 520 23 524
rect 277 520 280 524
rect 21 519 280 520
rect 21 515 23 519
rect 277 515 280 519
rect 21 514 280 515
rect 21 510 23 514
rect 277 510 280 514
rect 21 509 280 510
rect 21 505 23 509
rect 277 505 280 509
rect 21 504 280 505
rect 21 500 23 504
rect 277 500 280 504
rect 21 499 280 500
rect 21 495 23 499
rect 277 495 280 499
rect 21 494 280 495
rect 21 490 23 494
rect 277 490 280 494
rect 21 489 280 490
rect 21 485 23 489
rect 277 485 280 489
rect 21 484 280 485
rect 21 480 23 484
rect 277 480 280 484
rect 21 479 280 480
rect 21 475 23 479
rect 277 475 280 479
rect 21 474 280 475
rect 21 470 23 474
rect 277 470 280 474
rect 21 469 280 470
rect 21 465 23 469
rect 277 465 280 469
rect 21 464 280 465
rect 21 460 23 464
rect 277 460 280 464
rect 21 459 280 460
rect 21 455 23 459
rect 277 455 280 459
rect 21 454 280 455
rect 21 450 23 454
rect 277 450 280 454
rect 21 449 280 450
rect 21 445 23 449
rect 277 445 280 449
rect 21 444 280 445
rect 21 440 23 444
rect 277 440 280 444
rect 21 439 280 440
rect 21 435 23 439
rect 277 435 280 439
rect 21 433 280 435
rect 0 419 10 424
rect 102 424 198 433
rect 0 418 99 419
rect 0 414 2 418
rect 96 414 99 418
rect 0 413 99 414
rect 0 409 2 413
rect 96 409 99 413
rect 0 408 99 409
rect 0 404 2 408
rect 96 404 99 408
rect 0 403 99 404
rect 0 399 2 403
rect 96 399 99 403
rect 0 398 99 399
rect 0 394 2 398
rect 96 394 99 398
rect 0 393 99 394
rect 0 389 2 393
rect 96 389 99 393
rect 0 388 99 389
rect 0 384 2 388
rect 96 384 99 388
rect 0 383 99 384
rect 0 379 2 383
rect 96 379 99 383
rect 0 378 99 379
rect 0 374 2 378
rect 96 374 99 378
rect 0 373 99 374
rect 0 369 2 373
rect 96 369 99 373
rect 0 368 99 369
rect 0 364 2 368
rect 96 364 99 368
rect 0 363 99 364
rect 0 359 2 363
rect 96 359 99 363
rect 0 358 99 359
rect 0 349 2 358
rect 96 349 99 358
rect 0 348 99 349
rect 0 344 2 348
rect 96 344 99 348
rect 102 340 140 424
rect 143 418 157 421
rect 143 413 157 414
rect 143 408 157 409
rect 143 403 157 404
rect 143 398 157 399
rect 143 393 157 394
rect 143 388 157 389
rect 143 383 157 384
rect 143 378 157 379
rect 143 373 157 374
rect 143 368 157 369
rect 143 363 157 364
rect 143 358 157 359
rect 143 353 157 354
rect 143 348 157 349
rect 160 340 198 424
rect 289 424 290 658
rect 299 424 300 658
rect 289 419 300 424
rect 201 418 300 419
rect 201 414 204 418
rect 298 414 300 418
rect 201 413 300 414
rect 201 409 204 413
rect 298 409 300 413
rect 201 408 300 409
rect 201 404 204 408
rect 298 404 300 408
rect 201 403 300 404
rect 201 399 204 403
rect 298 399 300 403
rect 201 398 300 399
rect 201 394 204 398
rect 298 394 300 398
rect 201 393 300 394
rect 201 389 204 393
rect 298 389 300 393
rect 201 388 300 389
rect 201 384 204 388
rect 298 384 300 388
rect 201 383 300 384
rect 201 379 204 383
rect 298 379 300 383
rect 201 378 300 379
rect 201 374 204 378
rect 298 374 300 378
rect 201 373 300 374
rect 201 369 204 373
rect 298 369 300 373
rect 201 368 300 369
rect 201 364 204 368
rect 298 364 300 368
rect 201 363 300 364
rect 201 359 204 363
rect 298 359 300 363
rect 201 358 300 359
rect 201 354 204 358
rect 298 354 300 358
rect 201 353 300 354
rect 201 349 204 353
rect 298 349 300 353
rect 201 348 300 349
rect 201 344 204 348
rect 298 344 300 348
rect 102 326 198 340
rect 0 322 3 326
rect 297 322 300 326
rect 0 321 300 322
rect 0 317 3 321
rect 297 317 300 321
rect 0 316 300 317
rect 0 312 3 316
rect 297 312 300 316
rect 0 311 300 312
rect 0 307 3 311
rect 297 307 300 311
rect 0 306 300 307
rect 0 302 3 306
rect 297 302 300 306
rect 0 301 300 302
rect 0 297 3 301
rect 297 297 300 301
rect 0 296 300 297
rect 0 292 3 296
rect 297 292 300 296
rect 0 291 300 292
rect 0 287 3 291
rect 297 287 300 291
rect 0 286 300 287
rect 0 282 3 286
rect 297 282 300 286
rect 0 281 300 282
rect 0 277 3 281
rect 297 277 300 281
rect 0 276 300 277
rect 0 272 3 276
rect 297 272 300 276
rect 0 271 300 272
rect 0 267 3 271
rect 297 267 300 271
rect 0 266 300 267
rect 0 262 3 266
rect 297 262 300 266
rect 0 261 300 262
rect 0 257 8 261
rect 292 257 300 261
rect 0 256 300 257
rect 0 3 2 256
rect 6 252 8 256
rect 292 252 294 256
rect 6 251 294 252
rect 6 8 8 251
rect 14 241 99 246
rect 14 237 19 241
rect 98 237 99 241
rect 14 233 99 237
rect 14 228 24 233
rect 14 29 19 228
rect 23 29 24 228
rect 28 229 39 233
rect 98 229 99 233
rect 28 227 99 229
rect 28 223 41 227
rect 95 223 99 227
rect 28 217 99 223
rect 28 43 32 217
rect 36 215 99 217
rect 36 196 39 215
rect 53 211 57 215
rect 96 211 99 215
rect 102 230 198 251
rect 102 208 142 230
rect 36 194 53 196
rect 36 175 39 194
rect 56 200 142 208
rect 157 208 198 230
rect 201 244 286 246
rect 201 235 202 244
rect 281 235 286 244
rect 201 233 286 235
rect 201 229 202 233
rect 261 229 277 233
rect 201 228 277 229
rect 201 227 272 228
rect 201 223 205 227
rect 259 223 272 227
rect 201 217 272 223
rect 201 215 264 217
rect 201 211 204 215
rect 243 211 247 215
rect 157 200 244 208
rect 120 196 180 200
rect 56 194 244 196
rect 120 190 180 194
rect 56 182 244 190
rect 261 196 264 215
rect 247 194 264 196
rect 53 175 57 179
rect 116 175 120 179
rect 36 167 120 175
rect 36 163 41 167
rect 36 161 120 163
rect 36 157 41 161
rect 36 149 120 157
rect 36 110 39 149
rect 53 145 57 149
rect 116 145 120 149
rect 123 142 177 182
rect 180 175 184 179
rect 243 175 247 179
rect 261 175 264 194
rect 180 167 264 175
rect 259 163 264 167
rect 180 161 264 163
rect 259 157 264 161
rect 180 149 264 157
rect 180 145 184 149
rect 243 145 247 149
rect 56 138 244 142
rect 56 134 142 138
rect 120 125 142 134
rect 56 120 142 125
rect 157 134 244 138
rect 157 125 180 134
rect 157 120 244 125
rect 56 117 244 120
rect 53 110 57 114
rect 116 110 120 114
rect 36 102 120 110
rect 36 98 41 102
rect 36 96 120 98
rect 36 92 41 96
rect 36 84 120 92
rect 36 45 39 84
rect 53 80 57 84
rect 116 80 120 84
rect 123 77 177 117
rect 180 110 184 114
rect 243 110 247 114
rect 261 110 264 149
rect 180 102 264 110
rect 259 98 264 102
rect 180 96 264 98
rect 259 92 264 96
rect 180 84 264 92
rect 180 80 184 84
rect 243 80 247 84
rect 56 70 244 77
rect 56 69 142 70
rect 120 60 142 69
rect 157 69 244 70
rect 56 52 142 60
rect 53 45 57 49
rect 96 45 99 49
rect 36 43 99 45
rect 28 37 99 43
rect 28 33 41 37
rect 95 33 99 37
rect 28 29 39 33
rect 98 29 99 33
rect 14 27 99 29
rect 14 23 19 27
rect 98 23 99 27
rect 14 22 99 23
rect 14 18 19 22
rect 98 18 99 22
rect 14 14 99 18
rect 102 28 142 52
rect 157 60 180 69
rect 157 52 244 60
rect 157 28 198 52
rect 6 7 99 8
rect 6 3 8 7
rect 92 3 99 7
rect 0 0 99 3
rect 102 0 198 28
rect 201 45 204 49
rect 243 45 247 49
rect 261 45 264 84
rect 201 43 264 45
rect 268 43 272 217
rect 201 37 272 43
rect 201 33 205 37
rect 259 33 272 37
rect 201 29 202 33
rect 261 29 272 33
rect 276 29 277 228
rect 281 29 286 233
rect 201 27 286 29
rect 201 23 202 27
rect 281 23 286 27
rect 201 22 286 23
rect 201 18 202 22
rect 281 18 286 22
rect 201 14 286 18
rect 292 8 294 251
rect 201 7 294 8
rect 201 3 203 7
rect 292 3 294 7
rect 298 3 300 256
rect 201 0 300 3
<< m2contact >>
rect 23 640 277 644
rect 23 630 277 634
rect 23 620 277 624
rect 23 610 277 614
rect 23 600 277 604
rect 23 590 277 594
rect 23 580 277 584
rect 23 570 277 574
rect 23 560 277 564
rect 23 550 277 554
rect 23 540 277 544
rect 23 530 277 534
rect 23 520 277 524
rect 23 510 277 514
rect 23 500 277 504
rect 23 490 277 494
rect 23 480 277 484
rect 23 470 277 474
rect 23 460 277 464
rect 23 450 277 454
rect 23 440 277 444
rect 2 414 96 418
rect 2 404 96 408
rect 2 394 96 398
rect 2 384 96 388
rect 2 374 96 378
rect 2 364 96 368
rect 2 349 96 358
rect 143 409 157 413
rect 143 399 157 403
rect 143 389 157 393
rect 143 379 157 383
rect 143 369 157 373
rect 143 359 157 363
rect 143 349 157 353
rect 204 409 298 413
rect 204 399 298 403
rect 204 389 298 393
rect 204 379 298 383
rect 204 369 298 373
rect 204 359 298 363
rect 204 349 298 353
rect 3 317 297 321
rect 3 307 297 311
rect 3 297 297 301
rect 3 287 297 291
rect 3 277 297 281
rect 3 267 297 271
rect 8 257 292 261
rect 19 29 23 228
rect 39 196 53 215
rect 57 211 96 215
rect 39 175 53 194
rect 145 223 154 227
rect 145 215 154 219
rect 145 207 154 211
rect 204 211 243 215
rect 247 196 261 215
rect 57 175 116 179
rect 39 110 53 149
rect 57 145 116 149
rect 184 175 243 179
rect 247 175 261 194
rect 184 145 243 149
rect 145 127 154 131
rect 57 110 116 114
rect 39 45 53 84
rect 57 80 116 84
rect 184 110 243 114
rect 247 110 261 149
rect 184 80 243 84
rect 57 45 96 49
rect 39 29 98 33
rect 19 18 98 22
rect 145 63 154 67
rect 145 55 154 59
rect 145 47 154 51
rect 145 39 154 43
rect 145 31 154 35
rect 204 45 243 49
rect 247 45 261 84
rect 202 29 261 33
rect 272 29 276 228
rect 202 18 281 22
<< metal2 >>
rect 20 997 280 1000
rect 20 743 23 997
rect 277 743 280 997
rect 20 740 280 743
rect 0 644 300 670
rect 0 640 23 644
rect 277 640 300 644
rect 0 634 300 640
rect 0 630 23 634
rect 277 630 300 634
rect 0 624 300 630
rect 0 620 23 624
rect 277 620 300 624
rect 0 614 300 620
rect 0 610 23 614
rect 277 610 300 614
rect 0 604 300 610
rect 0 600 23 604
rect 277 600 300 604
rect 0 594 300 600
rect 0 590 23 594
rect 277 590 300 594
rect 0 584 300 590
rect 0 580 23 584
rect 277 580 300 584
rect 0 574 300 580
rect 0 570 23 574
rect 277 570 300 574
rect 0 564 300 570
rect 0 560 23 564
rect 277 560 300 564
rect 0 554 300 560
rect 0 550 23 554
rect 277 550 300 554
rect 0 544 300 550
rect 0 540 23 544
rect 277 540 300 544
rect 0 534 300 540
rect 0 530 23 534
rect 277 530 300 534
rect 0 524 300 530
rect 0 520 23 524
rect 277 520 300 524
rect 0 514 300 520
rect 0 510 23 514
rect 277 510 300 514
rect 0 504 300 510
rect 0 500 23 504
rect 277 500 300 504
rect 0 494 300 500
rect 0 490 23 494
rect 277 490 300 494
rect 0 484 300 490
rect 0 480 23 484
rect 277 480 300 484
rect 0 474 300 480
rect 0 470 23 474
rect 277 470 300 474
rect 0 464 300 470
rect 0 460 23 464
rect 277 460 300 464
rect 0 454 300 460
rect 0 450 23 454
rect 277 450 300 454
rect 0 444 300 450
rect 0 440 23 444
rect 277 440 300 444
rect 0 418 300 424
rect 0 414 2 418
rect 96 414 300 418
rect 0 413 300 414
rect 0 409 143 413
rect 157 409 204 413
rect 298 409 300 413
rect 0 408 300 409
rect 0 404 2 408
rect 96 404 300 408
rect 0 403 300 404
rect 0 399 143 403
rect 157 399 204 403
rect 298 399 300 403
rect 0 398 300 399
rect 0 394 2 398
rect 96 394 300 398
rect 0 393 300 394
rect 0 389 143 393
rect 157 389 204 393
rect 298 389 300 393
rect 0 388 300 389
rect 0 384 2 388
rect 96 384 300 388
rect 0 383 300 384
rect 0 379 143 383
rect 157 379 204 383
rect 298 379 300 383
rect 0 378 300 379
rect 0 374 2 378
rect 96 374 300 378
rect 0 373 300 374
rect 0 369 143 373
rect 157 369 204 373
rect 298 369 300 373
rect 0 368 300 369
rect 0 364 2 368
rect 96 364 300 368
rect 0 363 300 364
rect 0 359 143 363
rect 157 359 204 363
rect 298 359 300 363
rect 0 358 300 359
rect 0 349 2 358
rect 96 353 300 358
rect 96 349 143 353
rect 157 349 204 353
rect 298 349 300 353
rect 0 344 300 349
rect 0 321 300 326
rect 0 317 3 321
rect 297 317 300 321
rect 0 311 300 317
rect 0 307 3 311
rect 297 307 300 311
rect 0 301 300 307
rect 0 297 3 301
rect 297 297 300 301
rect 0 291 300 297
rect 0 287 3 291
rect 297 287 300 291
rect 0 281 300 287
rect 0 277 3 281
rect 297 277 300 281
rect 0 271 300 277
rect 0 267 3 271
rect 297 267 300 271
rect 0 261 300 267
rect 0 257 8 261
rect 292 257 300 261
rect 0 246 300 257
rect 0 228 300 230
rect 0 29 19 228
rect 23 227 272 228
rect 23 223 145 227
rect 154 223 272 227
rect 23 219 272 223
rect 23 215 145 219
rect 154 215 272 219
rect 23 196 39 215
rect 53 211 57 215
rect 96 211 204 215
rect 243 211 247 215
rect 53 207 145 211
rect 154 207 247 211
rect 53 196 247 207
rect 261 196 272 215
rect 23 194 272 196
rect 23 175 39 194
rect 53 179 247 194
rect 53 175 57 179
rect 116 175 184 179
rect 243 175 247 179
rect 261 175 272 194
rect 23 149 272 175
rect 23 110 39 149
rect 53 145 57 149
rect 116 145 184 149
rect 243 145 247 149
rect 53 131 247 145
rect 53 127 145 131
rect 154 127 247 131
rect 53 114 247 127
rect 53 110 57 114
rect 116 110 184 114
rect 243 110 247 114
rect 261 110 272 149
rect 23 84 272 110
rect 23 45 39 84
rect 53 80 57 84
rect 116 80 184 84
rect 243 80 247 84
rect 53 67 247 80
rect 53 63 145 67
rect 154 63 247 67
rect 53 59 247 63
rect 53 55 145 59
rect 154 55 247 59
rect 53 51 247 55
rect 53 49 145 51
rect 53 45 57 49
rect 96 47 145 49
rect 154 49 247 51
rect 154 47 204 49
rect 96 45 204 47
rect 243 45 247 49
rect 261 45 272 84
rect 23 43 272 45
rect 23 39 145 43
rect 154 39 272 43
rect 23 35 272 39
rect 23 33 145 35
rect 23 29 39 33
rect 98 31 145 33
rect 154 33 272 35
rect 154 31 202 33
rect 98 29 202 31
rect 261 29 272 33
rect 276 29 300 228
rect 0 22 300 29
rect 0 18 19 22
rect 98 18 202 22
rect 281 18 300 22
rect 0 7 300 18
rect 0 0 98 7
rect 202 0 300 7
<< pad >>
rect 23 743 277 997
<< m1p >>
rect 102 0 198 4
<< m3p >>
rect 130 855 143 868
<< labels >>
rlabel m3p 136 861 136 861 1 YPAD
rlabel m1p 150 0 150 0 8 vdd
<< end >>

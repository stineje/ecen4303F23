magic
tech  scmos
timestamp 777777777
<< poly >>
rect 180 553 181 554
rect 181 553 182 554
rect 182 553 183 554
rect 183 553 184 554
rect 184 553 185 554
rect 185 553 186 554
rect 186 553 187 554
rect 187 553 188 554
rect 188 553 189 554
rect 189 553 190 554
rect 176 552 177 553
rect 177 552 178 553
rect 178 552 179 553
rect 179 552 180 553
rect 180 552 181 553
rect 181 552 182 553
rect 182 552 183 553
rect 183 552 184 553
rect 184 552 185 553
rect 185 552 186 553
rect 186 552 187 553
rect 187 552 188 553
rect 188 552 189 553
rect 189 552 190 553
rect 190 552 191 553
rect 191 552 192 553
rect 192 552 193 553
rect 193 552 194 553
rect 174 551 175 552
rect 175 551 176 552
rect 176 551 177 552
rect 177 551 178 552
rect 178 551 179 552
rect 179 551 180 552
rect 180 551 181 552
rect 181 551 182 552
rect 182 551 183 552
rect 183 551 184 552
rect 184 551 185 552
rect 185 551 186 552
rect 186 551 187 552
rect 187 551 188 552
rect 188 551 189 552
rect 189 551 190 552
rect 190 551 191 552
rect 191 551 192 552
rect 192 551 193 552
rect 193 551 194 552
rect 194 551 195 552
rect 195 551 196 552
rect 196 551 197 552
rect 172 550 173 551
rect 173 550 174 551
rect 174 550 175 551
rect 175 550 176 551
rect 176 550 177 551
rect 177 550 178 551
rect 178 550 179 551
rect 179 550 180 551
rect 180 550 181 551
rect 181 550 182 551
rect 182 550 183 551
rect 183 550 184 551
rect 184 550 185 551
rect 185 550 186 551
rect 186 550 187 551
rect 187 550 188 551
rect 188 550 189 551
rect 189 550 190 551
rect 190 550 191 551
rect 191 550 192 551
rect 192 550 193 551
rect 193 550 194 551
rect 194 550 195 551
rect 195 550 196 551
rect 196 550 197 551
rect 197 550 198 551
rect 198 550 199 551
rect 199 550 200 551
rect 170 549 171 550
rect 171 549 172 550
rect 172 549 173 550
rect 173 549 174 550
rect 174 549 175 550
rect 175 549 176 550
rect 176 549 177 550
rect 177 549 178 550
rect 178 549 179 550
rect 179 549 180 550
rect 180 549 181 550
rect 181 549 182 550
rect 182 549 183 550
rect 183 549 184 550
rect 184 549 185 550
rect 185 549 186 550
rect 186 549 187 550
rect 187 549 188 550
rect 188 549 189 550
rect 189 549 190 550
rect 190 549 191 550
rect 191 549 192 550
rect 192 549 193 550
rect 193 549 194 550
rect 194 549 195 550
rect 195 549 196 550
rect 196 549 197 550
rect 197 549 198 550
rect 198 549 199 550
rect 199 549 200 550
rect 200 549 201 550
rect 201 549 202 550
rect 202 549 203 550
rect 169 548 170 549
rect 170 548 171 549
rect 171 548 172 549
rect 172 548 173 549
rect 173 548 174 549
rect 174 548 175 549
rect 175 548 176 549
rect 176 548 177 549
rect 177 548 178 549
rect 178 548 179 549
rect 179 548 180 549
rect 180 548 181 549
rect 181 548 182 549
rect 182 548 183 549
rect 183 548 184 549
rect 184 548 185 549
rect 185 548 186 549
rect 186 548 187 549
rect 187 548 188 549
rect 188 548 189 549
rect 189 548 190 549
rect 190 548 191 549
rect 191 548 192 549
rect 192 548 193 549
rect 193 548 194 549
rect 194 548 195 549
rect 195 548 196 549
rect 196 548 197 549
rect 197 548 198 549
rect 198 548 199 549
rect 199 548 200 549
rect 200 548 201 549
rect 201 548 202 549
rect 202 548 203 549
rect 203 548 204 549
rect 204 548 205 549
rect 205 548 206 549
rect 168 547 169 548
rect 169 547 170 548
rect 170 547 171 548
rect 171 547 172 548
rect 172 547 173 548
rect 173 547 174 548
rect 174 547 175 548
rect 175 547 176 548
rect 176 547 177 548
rect 177 547 178 548
rect 178 547 179 548
rect 179 547 180 548
rect 180 547 181 548
rect 181 547 182 548
rect 182 547 183 548
rect 183 547 184 548
rect 184 547 185 548
rect 185 547 186 548
rect 186 547 187 548
rect 187 547 188 548
rect 188 547 189 548
rect 189 547 190 548
rect 190 547 191 548
rect 191 547 192 548
rect 192 547 193 548
rect 193 547 194 548
rect 194 547 195 548
rect 195 547 196 548
rect 196 547 197 548
rect 197 547 198 548
rect 198 547 199 548
rect 199 547 200 548
rect 200 547 201 548
rect 201 547 202 548
rect 202 547 203 548
rect 203 547 204 548
rect 204 547 205 548
rect 205 547 206 548
rect 206 547 207 548
rect 207 547 208 548
rect 167 546 168 547
rect 168 546 169 547
rect 169 546 170 547
rect 170 546 171 547
rect 171 546 172 547
rect 172 546 173 547
rect 173 546 174 547
rect 174 546 175 547
rect 175 546 176 547
rect 176 546 177 547
rect 177 546 178 547
rect 178 546 179 547
rect 179 546 180 547
rect 180 546 181 547
rect 181 546 182 547
rect 182 546 183 547
rect 183 546 184 547
rect 184 546 185 547
rect 185 546 186 547
rect 186 546 187 547
rect 187 546 188 547
rect 188 546 189 547
rect 189 546 190 547
rect 190 546 191 547
rect 191 546 192 547
rect 192 546 193 547
rect 193 546 194 547
rect 194 546 195 547
rect 195 546 196 547
rect 196 546 197 547
rect 197 546 198 547
rect 198 546 199 547
rect 199 546 200 547
rect 200 546 201 547
rect 201 546 202 547
rect 202 546 203 547
rect 203 546 204 547
rect 204 546 205 547
rect 205 546 206 547
rect 206 546 207 547
rect 207 546 208 547
rect 208 546 209 547
rect 209 546 210 547
rect 210 546 211 547
rect 166 545 167 546
rect 167 545 168 546
rect 168 545 169 546
rect 169 545 170 546
rect 170 545 171 546
rect 171 545 172 546
rect 172 545 173 546
rect 173 545 174 546
rect 174 545 175 546
rect 175 545 176 546
rect 176 545 177 546
rect 177 545 178 546
rect 178 545 179 546
rect 179 545 180 546
rect 180 545 181 546
rect 181 545 182 546
rect 182 545 183 546
rect 183 545 184 546
rect 184 545 185 546
rect 185 545 186 546
rect 186 545 187 546
rect 187 545 188 546
rect 188 545 189 546
rect 189 545 190 546
rect 190 545 191 546
rect 191 545 192 546
rect 192 545 193 546
rect 193 545 194 546
rect 194 545 195 546
rect 195 545 196 546
rect 196 545 197 546
rect 197 545 198 546
rect 198 545 199 546
rect 199 545 200 546
rect 200 545 201 546
rect 201 545 202 546
rect 202 545 203 546
rect 203 545 204 546
rect 204 545 205 546
rect 205 545 206 546
rect 206 545 207 546
rect 207 545 208 546
rect 208 545 209 546
rect 209 545 210 546
rect 210 545 211 546
rect 211 545 212 546
rect 212 545 213 546
rect 165 544 166 545
rect 166 544 167 545
rect 167 544 168 545
rect 168 544 169 545
rect 169 544 170 545
rect 170 544 171 545
rect 171 544 172 545
rect 172 544 173 545
rect 173 544 174 545
rect 174 544 175 545
rect 175 544 176 545
rect 176 544 177 545
rect 177 544 178 545
rect 178 544 179 545
rect 179 544 180 545
rect 191 544 192 545
rect 192 544 193 545
rect 193 544 194 545
rect 194 544 195 545
rect 195 544 196 545
rect 196 544 197 545
rect 197 544 198 545
rect 198 544 199 545
rect 199 544 200 545
rect 200 544 201 545
rect 201 544 202 545
rect 202 544 203 545
rect 203 544 204 545
rect 204 544 205 545
rect 205 544 206 545
rect 206 544 207 545
rect 207 544 208 545
rect 208 544 209 545
rect 209 544 210 545
rect 210 544 211 545
rect 211 544 212 545
rect 212 544 213 545
rect 213 544 214 545
rect 214 544 215 545
rect 215 544 216 545
rect 164 543 165 544
rect 165 543 166 544
rect 166 543 167 544
rect 167 543 168 544
rect 168 543 169 544
rect 169 543 170 544
rect 170 543 171 544
rect 171 543 172 544
rect 172 543 173 544
rect 173 543 174 544
rect 174 543 175 544
rect 175 543 176 544
rect 176 543 177 544
rect 177 543 178 544
rect 194 543 195 544
rect 195 543 196 544
rect 196 543 197 544
rect 197 543 198 544
rect 198 543 199 544
rect 199 543 200 544
rect 200 543 201 544
rect 201 543 202 544
rect 202 543 203 544
rect 203 543 204 544
rect 204 543 205 544
rect 205 543 206 544
rect 206 543 207 544
rect 207 543 208 544
rect 208 543 209 544
rect 209 543 210 544
rect 210 543 211 544
rect 211 543 212 544
rect 212 543 213 544
rect 213 543 214 544
rect 214 543 215 544
rect 215 543 216 544
rect 216 543 217 544
rect 217 543 218 544
rect 163 542 164 543
rect 164 542 165 543
rect 165 542 166 543
rect 166 542 167 543
rect 167 542 168 543
rect 168 542 169 543
rect 169 542 170 543
rect 170 542 171 543
rect 171 542 172 543
rect 172 542 173 543
rect 173 542 174 543
rect 174 542 175 543
rect 175 542 176 543
rect 197 542 198 543
rect 198 542 199 543
rect 199 542 200 543
rect 200 542 201 543
rect 201 542 202 543
rect 202 542 203 543
rect 203 542 204 543
rect 204 542 205 543
rect 205 542 206 543
rect 206 542 207 543
rect 207 542 208 543
rect 208 542 209 543
rect 209 542 210 543
rect 210 542 211 543
rect 211 542 212 543
rect 212 542 213 543
rect 213 542 214 543
rect 214 542 215 543
rect 215 542 216 543
rect 216 542 217 543
rect 217 542 218 543
rect 218 542 219 543
rect 219 542 220 543
rect 162 541 163 542
rect 163 541 164 542
rect 164 541 165 542
rect 165 541 166 542
rect 166 541 167 542
rect 167 541 168 542
rect 168 541 169 542
rect 169 541 170 542
rect 170 541 171 542
rect 171 541 172 542
rect 172 541 173 542
rect 173 541 174 542
rect 174 541 175 542
rect 200 541 201 542
rect 201 541 202 542
rect 202 541 203 542
rect 203 541 204 542
rect 204 541 205 542
rect 205 541 206 542
rect 206 541 207 542
rect 207 541 208 542
rect 208 541 209 542
rect 209 541 210 542
rect 210 541 211 542
rect 211 541 212 542
rect 212 541 213 542
rect 213 541 214 542
rect 214 541 215 542
rect 215 541 216 542
rect 216 541 217 542
rect 217 541 218 542
rect 218 541 219 542
rect 219 541 220 542
rect 220 541 221 542
rect 221 541 222 542
rect 222 541 223 542
rect 161 540 162 541
rect 162 540 163 541
rect 163 540 164 541
rect 164 540 165 541
rect 165 540 166 541
rect 166 540 167 541
rect 167 540 168 541
rect 168 540 169 541
rect 169 540 170 541
rect 170 540 171 541
rect 171 540 172 541
rect 172 540 173 541
rect 203 540 204 541
rect 204 540 205 541
rect 205 540 206 541
rect 206 540 207 541
rect 207 540 208 541
rect 208 540 209 541
rect 209 540 210 541
rect 210 540 211 541
rect 211 540 212 541
rect 212 540 213 541
rect 213 540 214 541
rect 214 540 215 541
rect 215 540 216 541
rect 216 540 217 541
rect 217 540 218 541
rect 218 540 219 541
rect 219 540 220 541
rect 220 540 221 541
rect 221 540 222 541
rect 222 540 223 541
rect 223 540 224 541
rect 224 540 225 541
rect 161 539 162 540
rect 162 539 163 540
rect 163 539 164 540
rect 164 539 165 540
rect 165 539 166 540
rect 166 539 167 540
rect 167 539 168 540
rect 168 539 169 540
rect 169 539 170 540
rect 170 539 171 540
rect 171 539 172 540
rect 206 539 207 540
rect 207 539 208 540
rect 208 539 209 540
rect 209 539 210 540
rect 210 539 211 540
rect 211 539 212 540
rect 212 539 213 540
rect 213 539 214 540
rect 214 539 215 540
rect 215 539 216 540
rect 216 539 217 540
rect 217 539 218 540
rect 218 539 219 540
rect 219 539 220 540
rect 220 539 221 540
rect 221 539 222 540
rect 222 539 223 540
rect 223 539 224 540
rect 224 539 225 540
rect 225 539 226 540
rect 226 539 227 540
rect 160 538 161 539
rect 161 538 162 539
rect 162 538 163 539
rect 163 538 164 539
rect 164 538 165 539
rect 165 538 166 539
rect 166 538 167 539
rect 167 538 168 539
rect 168 538 169 539
rect 169 538 170 539
rect 170 538 171 539
rect 208 538 209 539
rect 209 538 210 539
rect 210 538 211 539
rect 211 538 212 539
rect 212 538 213 539
rect 213 538 214 539
rect 214 538 215 539
rect 215 538 216 539
rect 216 538 217 539
rect 217 538 218 539
rect 218 538 219 539
rect 219 538 220 539
rect 220 538 221 539
rect 221 538 222 539
rect 222 538 223 539
rect 223 538 224 539
rect 224 538 225 539
rect 225 538 226 539
rect 226 538 227 539
rect 227 538 228 539
rect 228 538 229 539
rect 159 537 160 538
rect 160 537 161 538
rect 161 537 162 538
rect 162 537 163 538
rect 163 537 164 538
rect 164 537 165 538
rect 165 537 166 538
rect 166 537 167 538
rect 167 537 168 538
rect 168 537 169 538
rect 169 537 170 538
rect 211 537 212 538
rect 212 537 213 538
rect 213 537 214 538
rect 214 537 215 538
rect 215 537 216 538
rect 216 537 217 538
rect 217 537 218 538
rect 218 537 219 538
rect 219 537 220 538
rect 220 537 221 538
rect 221 537 222 538
rect 222 537 223 538
rect 223 537 224 538
rect 224 537 225 538
rect 225 537 226 538
rect 226 537 227 538
rect 227 537 228 538
rect 228 537 229 538
rect 229 537 230 538
rect 230 537 231 538
rect 158 536 159 537
rect 159 536 160 537
rect 160 536 161 537
rect 161 536 162 537
rect 162 536 163 537
rect 163 536 164 537
rect 164 536 165 537
rect 165 536 166 537
rect 166 536 167 537
rect 167 536 168 537
rect 168 536 169 537
rect 169 536 170 537
rect 213 536 214 537
rect 214 536 215 537
rect 215 536 216 537
rect 216 536 217 537
rect 217 536 218 537
rect 218 536 219 537
rect 219 536 220 537
rect 220 536 221 537
rect 221 536 222 537
rect 222 536 223 537
rect 223 536 224 537
rect 224 536 225 537
rect 225 536 226 537
rect 226 536 227 537
rect 227 536 228 537
rect 228 536 229 537
rect 229 536 230 537
rect 230 536 231 537
rect 231 536 232 537
rect 232 536 233 537
rect 158 535 159 536
rect 159 535 160 536
rect 160 535 161 536
rect 161 535 162 536
rect 162 535 163 536
rect 163 535 164 536
rect 164 535 165 536
rect 165 535 166 536
rect 166 535 167 536
rect 167 535 168 536
rect 168 535 169 536
rect 215 535 216 536
rect 216 535 217 536
rect 217 535 218 536
rect 218 535 219 536
rect 219 535 220 536
rect 220 535 221 536
rect 221 535 222 536
rect 222 535 223 536
rect 223 535 224 536
rect 224 535 225 536
rect 225 535 226 536
rect 226 535 227 536
rect 227 535 228 536
rect 228 535 229 536
rect 229 535 230 536
rect 230 535 231 536
rect 231 535 232 536
rect 232 535 233 536
rect 233 535 234 536
rect 234 535 235 536
rect 157 534 158 535
rect 158 534 159 535
rect 159 534 160 535
rect 160 534 161 535
rect 161 534 162 535
rect 162 534 163 535
rect 163 534 164 535
rect 164 534 165 535
rect 165 534 166 535
rect 166 534 167 535
rect 167 534 168 535
rect 218 534 219 535
rect 219 534 220 535
rect 220 534 221 535
rect 221 534 222 535
rect 222 534 223 535
rect 223 534 224 535
rect 224 534 225 535
rect 225 534 226 535
rect 226 534 227 535
rect 227 534 228 535
rect 228 534 229 535
rect 229 534 230 535
rect 230 534 231 535
rect 231 534 232 535
rect 232 534 233 535
rect 233 534 234 535
rect 234 534 235 535
rect 235 534 236 535
rect 236 534 237 535
rect 156 533 157 534
rect 157 533 158 534
rect 158 533 159 534
rect 159 533 160 534
rect 160 533 161 534
rect 161 533 162 534
rect 162 533 163 534
rect 163 533 164 534
rect 164 533 165 534
rect 165 533 166 534
rect 166 533 167 534
rect 220 533 221 534
rect 221 533 222 534
rect 222 533 223 534
rect 223 533 224 534
rect 224 533 225 534
rect 225 533 226 534
rect 226 533 227 534
rect 227 533 228 534
rect 228 533 229 534
rect 229 533 230 534
rect 230 533 231 534
rect 231 533 232 534
rect 232 533 233 534
rect 233 533 234 534
rect 234 533 235 534
rect 235 533 236 534
rect 236 533 237 534
rect 237 533 238 534
rect 156 532 157 533
rect 157 532 158 533
rect 158 532 159 533
rect 159 532 160 533
rect 160 532 161 533
rect 161 532 162 533
rect 162 532 163 533
rect 163 532 164 533
rect 164 532 165 533
rect 165 532 166 533
rect 166 532 167 533
rect 222 532 223 533
rect 223 532 224 533
rect 224 532 225 533
rect 225 532 226 533
rect 226 532 227 533
rect 227 532 228 533
rect 228 532 229 533
rect 229 532 230 533
rect 230 532 231 533
rect 231 532 232 533
rect 232 532 233 533
rect 233 532 234 533
rect 234 532 235 533
rect 235 532 236 533
rect 236 532 237 533
rect 237 532 238 533
rect 238 532 239 533
rect 239 532 240 533
rect 155 531 156 532
rect 156 531 157 532
rect 157 531 158 532
rect 158 531 159 532
rect 159 531 160 532
rect 160 531 161 532
rect 161 531 162 532
rect 162 531 163 532
rect 163 531 164 532
rect 164 531 165 532
rect 165 531 166 532
rect 224 531 225 532
rect 225 531 226 532
rect 226 531 227 532
rect 227 531 228 532
rect 228 531 229 532
rect 229 531 230 532
rect 230 531 231 532
rect 231 531 232 532
rect 232 531 233 532
rect 233 531 234 532
rect 234 531 235 532
rect 235 531 236 532
rect 236 531 237 532
rect 237 531 238 532
rect 238 531 239 532
rect 239 531 240 532
rect 240 531 241 532
rect 241 531 242 532
rect 151 530 152 531
rect 152 530 153 531
rect 153 530 154 531
rect 154 530 155 531
rect 155 530 156 531
rect 156 530 157 531
rect 157 530 158 531
rect 158 530 159 531
rect 159 530 160 531
rect 160 530 161 531
rect 161 530 162 531
rect 162 530 163 531
rect 163 530 164 531
rect 164 530 165 531
rect 226 530 227 531
rect 227 530 228 531
rect 228 530 229 531
rect 229 530 230 531
rect 230 530 231 531
rect 231 530 232 531
rect 232 530 233 531
rect 233 530 234 531
rect 234 530 235 531
rect 235 530 236 531
rect 236 530 237 531
rect 237 530 238 531
rect 238 530 239 531
rect 239 530 240 531
rect 240 530 241 531
rect 241 530 242 531
rect 242 530 243 531
rect 243 530 244 531
rect 147 529 148 530
rect 148 529 149 530
rect 149 529 150 530
rect 150 529 151 530
rect 151 529 152 530
rect 152 529 153 530
rect 153 529 154 530
rect 154 529 155 530
rect 155 529 156 530
rect 156 529 157 530
rect 157 529 158 530
rect 158 529 159 530
rect 159 529 160 530
rect 160 529 161 530
rect 161 529 162 530
rect 162 529 163 530
rect 163 529 164 530
rect 228 529 229 530
rect 229 529 230 530
rect 230 529 231 530
rect 231 529 232 530
rect 232 529 233 530
rect 233 529 234 530
rect 234 529 235 530
rect 235 529 236 530
rect 236 529 237 530
rect 237 529 238 530
rect 238 529 239 530
rect 239 529 240 530
rect 240 529 241 530
rect 241 529 242 530
rect 242 529 243 530
rect 243 529 244 530
rect 244 529 245 530
rect 245 529 246 530
rect 144 528 145 529
rect 145 528 146 529
rect 146 528 147 529
rect 147 528 148 529
rect 148 528 149 529
rect 149 528 150 529
rect 150 528 151 529
rect 151 528 152 529
rect 152 528 153 529
rect 153 528 154 529
rect 154 528 155 529
rect 155 528 156 529
rect 156 528 157 529
rect 157 528 158 529
rect 158 528 159 529
rect 159 528 160 529
rect 160 528 161 529
rect 161 528 162 529
rect 162 528 163 529
rect 163 528 164 529
rect 230 528 231 529
rect 231 528 232 529
rect 232 528 233 529
rect 233 528 234 529
rect 234 528 235 529
rect 235 528 236 529
rect 236 528 237 529
rect 237 528 238 529
rect 238 528 239 529
rect 239 528 240 529
rect 240 528 241 529
rect 241 528 242 529
rect 242 528 243 529
rect 243 528 244 529
rect 244 528 245 529
rect 245 528 246 529
rect 246 528 247 529
rect 247 528 248 529
rect 141 527 142 528
rect 142 527 143 528
rect 143 527 144 528
rect 144 527 145 528
rect 145 527 146 528
rect 146 527 147 528
rect 147 527 148 528
rect 148 527 149 528
rect 149 527 150 528
rect 150 527 151 528
rect 151 527 152 528
rect 152 527 153 528
rect 153 527 154 528
rect 154 527 155 528
rect 155 527 156 528
rect 156 527 157 528
rect 157 527 158 528
rect 158 527 159 528
rect 159 527 160 528
rect 160 527 161 528
rect 161 527 162 528
rect 162 527 163 528
rect 232 527 233 528
rect 233 527 234 528
rect 234 527 235 528
rect 235 527 236 528
rect 236 527 237 528
rect 237 527 238 528
rect 238 527 239 528
rect 239 527 240 528
rect 240 527 241 528
rect 241 527 242 528
rect 242 527 243 528
rect 243 527 244 528
rect 244 527 245 528
rect 245 527 246 528
rect 246 527 247 528
rect 247 527 248 528
rect 248 527 249 528
rect 139 526 140 527
rect 140 526 141 527
rect 141 526 142 527
rect 142 526 143 527
rect 143 526 144 527
rect 144 526 145 527
rect 145 526 146 527
rect 146 526 147 527
rect 147 526 148 527
rect 148 526 149 527
rect 149 526 150 527
rect 150 526 151 527
rect 151 526 152 527
rect 152 526 153 527
rect 153 526 154 527
rect 154 526 155 527
rect 155 526 156 527
rect 156 526 157 527
rect 157 526 158 527
rect 158 526 159 527
rect 159 526 160 527
rect 160 526 161 527
rect 161 526 162 527
rect 234 526 235 527
rect 235 526 236 527
rect 236 526 237 527
rect 237 526 238 527
rect 238 526 239 527
rect 239 526 240 527
rect 240 526 241 527
rect 241 526 242 527
rect 242 526 243 527
rect 243 526 244 527
rect 244 526 245 527
rect 245 526 246 527
rect 246 526 247 527
rect 247 526 248 527
rect 248 526 249 527
rect 249 526 250 527
rect 250 526 251 527
rect 138 525 139 526
rect 139 525 140 526
rect 140 525 141 526
rect 141 525 142 526
rect 142 525 143 526
rect 143 525 144 526
rect 144 525 145 526
rect 145 525 146 526
rect 146 525 147 526
rect 147 525 148 526
rect 148 525 149 526
rect 149 525 150 526
rect 150 525 151 526
rect 151 525 152 526
rect 152 525 153 526
rect 153 525 154 526
rect 154 525 155 526
rect 155 525 156 526
rect 156 525 157 526
rect 157 525 158 526
rect 158 525 159 526
rect 159 525 160 526
rect 160 525 161 526
rect 161 525 162 526
rect 187 525 188 526
rect 236 525 237 526
rect 237 525 238 526
rect 238 525 239 526
rect 239 525 240 526
rect 240 525 241 526
rect 241 525 242 526
rect 242 525 243 526
rect 243 525 244 526
rect 244 525 245 526
rect 245 525 246 526
rect 246 525 247 526
rect 247 525 248 526
rect 248 525 249 526
rect 249 525 250 526
rect 250 525 251 526
rect 251 525 252 526
rect 252 525 253 526
rect 136 524 137 525
rect 137 524 138 525
rect 138 524 139 525
rect 139 524 140 525
rect 140 524 141 525
rect 141 524 142 525
rect 142 524 143 525
rect 143 524 144 525
rect 144 524 145 525
rect 145 524 146 525
rect 146 524 147 525
rect 147 524 148 525
rect 148 524 149 525
rect 149 524 150 525
rect 150 524 151 525
rect 151 524 152 525
rect 152 524 153 525
rect 153 524 154 525
rect 154 524 155 525
rect 155 524 156 525
rect 156 524 157 525
rect 157 524 158 525
rect 158 524 159 525
rect 159 524 160 525
rect 160 524 161 525
rect 187 524 188 525
rect 188 524 189 525
rect 237 524 238 525
rect 238 524 239 525
rect 239 524 240 525
rect 240 524 241 525
rect 241 524 242 525
rect 242 524 243 525
rect 243 524 244 525
rect 244 524 245 525
rect 245 524 246 525
rect 246 524 247 525
rect 247 524 248 525
rect 248 524 249 525
rect 249 524 250 525
rect 250 524 251 525
rect 251 524 252 525
rect 252 524 253 525
rect 253 524 254 525
rect 135 523 136 524
rect 136 523 137 524
rect 137 523 138 524
rect 138 523 139 524
rect 139 523 140 524
rect 140 523 141 524
rect 141 523 142 524
rect 142 523 143 524
rect 143 523 144 524
rect 144 523 145 524
rect 145 523 146 524
rect 146 523 147 524
rect 147 523 148 524
rect 148 523 149 524
rect 149 523 150 524
rect 150 523 151 524
rect 151 523 152 524
rect 152 523 153 524
rect 153 523 154 524
rect 154 523 155 524
rect 155 523 156 524
rect 156 523 157 524
rect 157 523 158 524
rect 158 523 159 524
rect 159 523 160 524
rect 160 523 161 524
rect 188 523 189 524
rect 189 523 190 524
rect 239 523 240 524
rect 240 523 241 524
rect 241 523 242 524
rect 242 523 243 524
rect 243 523 244 524
rect 244 523 245 524
rect 245 523 246 524
rect 246 523 247 524
rect 247 523 248 524
rect 248 523 249 524
rect 249 523 250 524
rect 250 523 251 524
rect 251 523 252 524
rect 252 523 253 524
rect 253 523 254 524
rect 254 523 255 524
rect 255 523 256 524
rect 134 522 135 523
rect 135 522 136 523
rect 136 522 137 523
rect 137 522 138 523
rect 138 522 139 523
rect 139 522 140 523
rect 140 522 141 523
rect 141 522 142 523
rect 142 522 143 523
rect 143 522 144 523
rect 144 522 145 523
rect 145 522 146 523
rect 146 522 147 523
rect 147 522 148 523
rect 148 522 149 523
rect 149 522 150 523
rect 150 522 151 523
rect 151 522 152 523
rect 152 522 153 523
rect 153 522 154 523
rect 154 522 155 523
rect 155 522 156 523
rect 156 522 157 523
rect 157 522 158 523
rect 158 522 159 523
rect 159 522 160 523
rect 189 522 190 523
rect 190 522 191 523
rect 241 522 242 523
rect 242 522 243 523
rect 243 522 244 523
rect 244 522 245 523
rect 245 522 246 523
rect 246 522 247 523
rect 247 522 248 523
rect 248 522 249 523
rect 249 522 250 523
rect 250 522 251 523
rect 251 522 252 523
rect 252 522 253 523
rect 253 522 254 523
rect 254 522 255 523
rect 255 522 256 523
rect 256 522 257 523
rect 257 522 258 523
rect 133 521 134 522
rect 134 521 135 522
rect 135 521 136 522
rect 136 521 137 522
rect 137 521 138 522
rect 138 521 139 522
rect 139 521 140 522
rect 140 521 141 522
rect 141 521 142 522
rect 142 521 143 522
rect 143 521 144 522
rect 144 521 145 522
rect 145 521 146 522
rect 146 521 147 522
rect 147 521 148 522
rect 148 521 149 522
rect 149 521 150 522
rect 150 521 151 522
rect 151 521 152 522
rect 152 521 153 522
rect 153 521 154 522
rect 154 521 155 522
rect 155 521 156 522
rect 156 521 157 522
rect 157 521 158 522
rect 158 521 159 522
rect 190 521 191 522
rect 191 521 192 522
rect 243 521 244 522
rect 244 521 245 522
rect 245 521 246 522
rect 246 521 247 522
rect 247 521 248 522
rect 248 521 249 522
rect 249 521 250 522
rect 250 521 251 522
rect 251 521 252 522
rect 252 521 253 522
rect 253 521 254 522
rect 254 521 255 522
rect 255 521 256 522
rect 256 521 257 522
rect 257 521 258 522
rect 258 521 259 522
rect 132 520 133 521
rect 133 520 134 521
rect 134 520 135 521
rect 135 520 136 521
rect 136 520 137 521
rect 137 520 138 521
rect 138 520 139 521
rect 139 520 140 521
rect 140 520 141 521
rect 141 520 142 521
rect 142 520 143 521
rect 143 520 144 521
rect 144 520 145 521
rect 145 520 146 521
rect 146 520 147 521
rect 147 520 148 521
rect 151 520 152 521
rect 152 520 153 521
rect 153 520 154 521
rect 154 520 155 521
rect 155 520 156 521
rect 156 520 157 521
rect 157 520 158 521
rect 158 520 159 521
rect 190 520 191 521
rect 191 520 192 521
rect 192 520 193 521
rect 245 520 246 521
rect 246 520 247 521
rect 247 520 248 521
rect 248 520 249 521
rect 249 520 250 521
rect 250 520 251 521
rect 251 520 252 521
rect 252 520 253 521
rect 253 520 254 521
rect 254 520 255 521
rect 255 520 256 521
rect 256 520 257 521
rect 257 520 258 521
rect 258 520 259 521
rect 259 520 260 521
rect 260 520 261 521
rect 132 519 133 520
rect 133 519 134 520
rect 134 519 135 520
rect 135 519 136 520
rect 136 519 137 520
rect 137 519 138 520
rect 138 519 139 520
rect 139 519 140 520
rect 140 519 141 520
rect 141 519 142 520
rect 142 519 143 520
rect 143 519 144 520
rect 144 519 145 520
rect 151 519 152 520
rect 152 519 153 520
rect 153 519 154 520
rect 154 519 155 520
rect 155 519 156 520
rect 156 519 157 520
rect 157 519 158 520
rect 191 519 192 520
rect 192 519 193 520
rect 193 519 194 520
rect 194 519 195 520
rect 246 519 247 520
rect 247 519 248 520
rect 248 519 249 520
rect 249 519 250 520
rect 250 519 251 520
rect 251 519 252 520
rect 252 519 253 520
rect 253 519 254 520
rect 254 519 255 520
rect 255 519 256 520
rect 256 519 257 520
rect 257 519 258 520
rect 258 519 259 520
rect 259 519 260 520
rect 260 519 261 520
rect 261 519 262 520
rect 262 519 263 520
rect 131 518 132 519
rect 132 518 133 519
rect 133 518 134 519
rect 134 518 135 519
rect 135 518 136 519
rect 136 518 137 519
rect 137 518 138 519
rect 138 518 139 519
rect 139 518 140 519
rect 140 518 141 519
rect 141 518 142 519
rect 142 518 143 519
rect 150 518 151 519
rect 151 518 152 519
rect 152 518 153 519
rect 153 518 154 519
rect 154 518 155 519
rect 155 518 156 519
rect 156 518 157 519
rect 157 518 158 519
rect 192 518 193 519
rect 193 518 194 519
rect 194 518 195 519
rect 195 518 196 519
rect 248 518 249 519
rect 249 518 250 519
rect 250 518 251 519
rect 251 518 252 519
rect 252 518 253 519
rect 253 518 254 519
rect 254 518 255 519
rect 255 518 256 519
rect 256 518 257 519
rect 257 518 258 519
rect 258 518 259 519
rect 259 518 260 519
rect 260 518 261 519
rect 261 518 262 519
rect 262 518 263 519
rect 263 518 264 519
rect 130 517 131 518
rect 131 517 132 518
rect 132 517 133 518
rect 133 517 134 518
rect 134 517 135 518
rect 135 517 136 518
rect 136 517 137 518
rect 137 517 138 518
rect 138 517 139 518
rect 139 517 140 518
rect 140 517 141 518
rect 141 517 142 518
rect 149 517 150 518
rect 150 517 151 518
rect 151 517 152 518
rect 152 517 153 518
rect 153 517 154 518
rect 154 517 155 518
rect 155 517 156 518
rect 156 517 157 518
rect 192 517 193 518
rect 193 517 194 518
rect 194 517 195 518
rect 195 517 196 518
rect 196 517 197 518
rect 250 517 251 518
rect 251 517 252 518
rect 252 517 253 518
rect 253 517 254 518
rect 254 517 255 518
rect 255 517 256 518
rect 256 517 257 518
rect 257 517 258 518
rect 258 517 259 518
rect 259 517 260 518
rect 260 517 261 518
rect 261 517 262 518
rect 262 517 263 518
rect 263 517 264 518
rect 264 517 265 518
rect 265 517 266 518
rect 130 516 131 517
rect 131 516 132 517
rect 132 516 133 517
rect 133 516 134 517
rect 134 516 135 517
rect 135 516 136 517
rect 136 516 137 517
rect 137 516 138 517
rect 138 516 139 517
rect 139 516 140 517
rect 140 516 141 517
rect 149 516 150 517
rect 150 516 151 517
rect 151 516 152 517
rect 152 516 153 517
rect 153 516 154 517
rect 154 516 155 517
rect 155 516 156 517
rect 193 516 194 517
rect 194 516 195 517
rect 195 516 196 517
rect 196 516 197 517
rect 197 516 198 517
rect 252 516 253 517
rect 253 516 254 517
rect 254 516 255 517
rect 255 516 256 517
rect 256 516 257 517
rect 257 516 258 517
rect 258 516 259 517
rect 259 516 260 517
rect 260 516 261 517
rect 261 516 262 517
rect 262 516 263 517
rect 263 516 264 517
rect 264 516 265 517
rect 265 516 266 517
rect 266 516 267 517
rect 267 516 268 517
rect 129 515 130 516
rect 130 515 131 516
rect 131 515 132 516
rect 132 515 133 516
rect 133 515 134 516
rect 134 515 135 516
rect 135 515 136 516
rect 136 515 137 516
rect 137 515 138 516
rect 138 515 139 516
rect 139 515 140 516
rect 148 515 149 516
rect 149 515 150 516
rect 150 515 151 516
rect 151 515 152 516
rect 152 515 153 516
rect 153 515 154 516
rect 154 515 155 516
rect 155 515 156 516
rect 194 515 195 516
rect 195 515 196 516
rect 196 515 197 516
rect 197 515 198 516
rect 198 515 199 516
rect 253 515 254 516
rect 254 515 255 516
rect 255 515 256 516
rect 256 515 257 516
rect 257 515 258 516
rect 258 515 259 516
rect 259 515 260 516
rect 260 515 261 516
rect 261 515 262 516
rect 262 515 263 516
rect 263 515 264 516
rect 264 515 265 516
rect 265 515 266 516
rect 266 515 267 516
rect 267 515 268 516
rect 268 515 269 516
rect 129 514 130 515
rect 130 514 131 515
rect 131 514 132 515
rect 132 514 133 515
rect 133 514 134 515
rect 134 514 135 515
rect 135 514 136 515
rect 136 514 137 515
rect 137 514 138 515
rect 138 514 139 515
rect 147 514 148 515
rect 148 514 149 515
rect 149 514 150 515
rect 150 514 151 515
rect 151 514 152 515
rect 152 514 153 515
rect 153 514 154 515
rect 154 514 155 515
rect 195 514 196 515
rect 196 514 197 515
rect 197 514 198 515
rect 198 514 199 515
rect 199 514 200 515
rect 255 514 256 515
rect 256 514 257 515
rect 257 514 258 515
rect 258 514 259 515
rect 259 514 260 515
rect 260 514 261 515
rect 261 514 262 515
rect 262 514 263 515
rect 263 514 264 515
rect 264 514 265 515
rect 265 514 266 515
rect 266 514 267 515
rect 267 514 268 515
rect 268 514 269 515
rect 269 514 270 515
rect 270 514 271 515
rect 129 513 130 514
rect 130 513 131 514
rect 131 513 132 514
rect 132 513 133 514
rect 133 513 134 514
rect 134 513 135 514
rect 135 513 136 514
rect 136 513 137 514
rect 137 513 138 514
rect 145 513 146 514
rect 146 513 147 514
rect 147 513 148 514
rect 148 513 149 514
rect 149 513 150 514
rect 150 513 151 514
rect 151 513 152 514
rect 152 513 153 514
rect 153 513 154 514
rect 195 513 196 514
rect 196 513 197 514
rect 197 513 198 514
rect 198 513 199 514
rect 199 513 200 514
rect 200 513 201 514
rect 201 513 202 514
rect 225 513 226 514
rect 257 513 258 514
rect 258 513 259 514
rect 259 513 260 514
rect 260 513 261 514
rect 261 513 262 514
rect 262 513 263 514
rect 263 513 264 514
rect 264 513 265 514
rect 265 513 266 514
rect 266 513 267 514
rect 267 513 268 514
rect 268 513 269 514
rect 269 513 270 514
rect 270 513 271 514
rect 271 513 272 514
rect 128 512 129 513
rect 129 512 130 513
rect 130 512 131 513
rect 131 512 132 513
rect 132 512 133 513
rect 133 512 134 513
rect 134 512 135 513
rect 135 512 136 513
rect 136 512 137 513
rect 137 512 138 513
rect 146 512 147 513
rect 147 512 148 513
rect 148 512 149 513
rect 149 512 150 513
rect 150 512 151 513
rect 151 512 152 513
rect 196 512 197 513
rect 197 512 198 513
rect 198 512 199 513
rect 199 512 200 513
rect 200 512 201 513
rect 201 512 202 513
rect 202 512 203 513
rect 225 512 226 513
rect 226 512 227 513
rect 258 512 259 513
rect 259 512 260 513
rect 260 512 261 513
rect 261 512 262 513
rect 262 512 263 513
rect 263 512 264 513
rect 264 512 265 513
rect 265 512 266 513
rect 266 512 267 513
rect 267 512 268 513
rect 268 512 269 513
rect 269 512 270 513
rect 270 512 271 513
rect 271 512 272 513
rect 272 512 273 513
rect 273 512 274 513
rect 128 511 129 512
rect 129 511 130 512
rect 130 511 131 512
rect 131 511 132 512
rect 132 511 133 512
rect 133 511 134 512
rect 134 511 135 512
rect 135 511 136 512
rect 136 511 137 512
rect 197 511 198 512
rect 198 511 199 512
rect 199 511 200 512
rect 200 511 201 512
rect 201 511 202 512
rect 202 511 203 512
rect 203 511 204 512
rect 225 511 226 512
rect 226 511 227 512
rect 227 511 228 512
rect 260 511 261 512
rect 261 511 262 512
rect 262 511 263 512
rect 263 511 264 512
rect 264 511 265 512
rect 265 511 266 512
rect 266 511 267 512
rect 267 511 268 512
rect 268 511 269 512
rect 269 511 270 512
rect 270 511 271 512
rect 271 511 272 512
rect 272 511 273 512
rect 273 511 274 512
rect 274 511 275 512
rect 275 511 276 512
rect 321 511 322 512
rect 322 511 323 512
rect 323 511 324 512
rect 324 511 325 512
rect 325 511 326 512
rect 326 511 327 512
rect 327 511 328 512
rect 328 511 329 512
rect 329 511 330 512
rect 330 511 331 512
rect 331 511 332 512
rect 332 511 333 512
rect 333 511 334 512
rect 334 511 335 512
rect 128 510 129 511
rect 129 510 130 511
rect 130 510 131 511
rect 131 510 132 511
rect 132 510 133 511
rect 133 510 134 511
rect 134 510 135 511
rect 135 510 136 511
rect 136 510 137 511
rect 197 510 198 511
rect 198 510 199 511
rect 199 510 200 511
rect 200 510 201 511
rect 201 510 202 511
rect 202 510 203 511
rect 203 510 204 511
rect 204 510 205 511
rect 226 510 227 511
rect 227 510 228 511
rect 228 510 229 511
rect 261 510 262 511
rect 262 510 263 511
rect 263 510 264 511
rect 264 510 265 511
rect 265 510 266 511
rect 266 510 267 511
rect 267 510 268 511
rect 268 510 269 511
rect 269 510 270 511
rect 270 510 271 511
rect 271 510 272 511
rect 272 510 273 511
rect 273 510 274 511
rect 274 510 275 511
rect 275 510 276 511
rect 276 510 277 511
rect 311 510 312 511
rect 312 510 313 511
rect 313 510 314 511
rect 314 510 315 511
rect 315 510 316 511
rect 316 510 317 511
rect 317 510 318 511
rect 318 510 319 511
rect 319 510 320 511
rect 320 510 321 511
rect 321 510 322 511
rect 322 510 323 511
rect 323 510 324 511
rect 324 510 325 511
rect 325 510 326 511
rect 326 510 327 511
rect 327 510 328 511
rect 328 510 329 511
rect 329 510 330 511
rect 330 510 331 511
rect 331 510 332 511
rect 332 510 333 511
rect 333 510 334 511
rect 334 510 335 511
rect 335 510 336 511
rect 336 510 337 511
rect 337 510 338 511
rect 338 510 339 511
rect 339 510 340 511
rect 340 510 341 511
rect 341 510 342 511
rect 342 510 343 511
rect 343 510 344 511
rect 128 509 129 510
rect 129 509 130 510
rect 130 509 131 510
rect 131 509 132 510
rect 132 509 133 510
rect 133 509 134 510
rect 134 509 135 510
rect 135 509 136 510
rect 136 509 137 510
rect 198 509 199 510
rect 199 509 200 510
rect 200 509 201 510
rect 201 509 202 510
rect 202 509 203 510
rect 203 509 204 510
rect 204 509 205 510
rect 205 509 206 510
rect 206 509 207 510
rect 226 509 227 510
rect 227 509 228 510
rect 228 509 229 510
rect 229 509 230 510
rect 230 509 231 510
rect 263 509 264 510
rect 264 509 265 510
rect 265 509 266 510
rect 266 509 267 510
rect 267 509 268 510
rect 268 509 269 510
rect 269 509 270 510
rect 270 509 271 510
rect 271 509 272 510
rect 272 509 273 510
rect 273 509 274 510
rect 274 509 275 510
rect 275 509 276 510
rect 276 509 277 510
rect 277 509 278 510
rect 278 509 279 510
rect 304 509 305 510
rect 305 509 306 510
rect 306 509 307 510
rect 307 509 308 510
rect 308 509 309 510
rect 309 509 310 510
rect 310 509 311 510
rect 311 509 312 510
rect 312 509 313 510
rect 313 509 314 510
rect 314 509 315 510
rect 315 509 316 510
rect 316 509 317 510
rect 317 509 318 510
rect 318 509 319 510
rect 319 509 320 510
rect 320 509 321 510
rect 321 509 322 510
rect 322 509 323 510
rect 323 509 324 510
rect 324 509 325 510
rect 325 509 326 510
rect 326 509 327 510
rect 327 509 328 510
rect 328 509 329 510
rect 329 509 330 510
rect 330 509 331 510
rect 331 509 332 510
rect 332 509 333 510
rect 333 509 334 510
rect 334 509 335 510
rect 335 509 336 510
rect 336 509 337 510
rect 337 509 338 510
rect 338 509 339 510
rect 339 509 340 510
rect 340 509 341 510
rect 341 509 342 510
rect 342 509 343 510
rect 343 509 344 510
rect 344 509 345 510
rect 345 509 346 510
rect 346 509 347 510
rect 347 509 348 510
rect 348 509 349 510
rect 349 509 350 510
rect 128 508 129 509
rect 129 508 130 509
rect 130 508 131 509
rect 131 508 132 509
rect 132 508 133 509
rect 133 508 134 509
rect 134 508 135 509
rect 135 508 136 509
rect 199 508 200 509
rect 200 508 201 509
rect 201 508 202 509
rect 202 508 203 509
rect 203 508 204 509
rect 204 508 205 509
rect 205 508 206 509
rect 206 508 207 509
rect 207 508 208 509
rect 226 508 227 509
rect 227 508 228 509
rect 228 508 229 509
rect 229 508 230 509
rect 230 508 231 509
rect 231 508 232 509
rect 265 508 266 509
rect 266 508 267 509
rect 267 508 268 509
rect 268 508 269 509
rect 269 508 270 509
rect 270 508 271 509
rect 271 508 272 509
rect 272 508 273 509
rect 273 508 274 509
rect 274 508 275 509
rect 275 508 276 509
rect 276 508 277 509
rect 277 508 278 509
rect 278 508 279 509
rect 279 508 280 509
rect 299 508 300 509
rect 300 508 301 509
rect 301 508 302 509
rect 302 508 303 509
rect 303 508 304 509
rect 304 508 305 509
rect 305 508 306 509
rect 306 508 307 509
rect 307 508 308 509
rect 308 508 309 509
rect 309 508 310 509
rect 310 508 311 509
rect 311 508 312 509
rect 312 508 313 509
rect 313 508 314 509
rect 314 508 315 509
rect 315 508 316 509
rect 316 508 317 509
rect 317 508 318 509
rect 318 508 319 509
rect 319 508 320 509
rect 320 508 321 509
rect 321 508 322 509
rect 322 508 323 509
rect 323 508 324 509
rect 324 508 325 509
rect 325 508 326 509
rect 326 508 327 509
rect 327 508 328 509
rect 328 508 329 509
rect 329 508 330 509
rect 330 508 331 509
rect 331 508 332 509
rect 332 508 333 509
rect 333 508 334 509
rect 334 508 335 509
rect 335 508 336 509
rect 336 508 337 509
rect 337 508 338 509
rect 338 508 339 509
rect 339 508 340 509
rect 340 508 341 509
rect 341 508 342 509
rect 342 508 343 509
rect 343 508 344 509
rect 344 508 345 509
rect 345 508 346 509
rect 346 508 347 509
rect 347 508 348 509
rect 348 508 349 509
rect 349 508 350 509
rect 350 508 351 509
rect 351 508 352 509
rect 352 508 353 509
rect 127 507 128 508
rect 128 507 129 508
rect 129 507 130 508
rect 130 507 131 508
rect 131 507 132 508
rect 132 507 133 508
rect 133 507 134 508
rect 134 507 135 508
rect 135 507 136 508
rect 199 507 200 508
rect 200 507 201 508
rect 201 507 202 508
rect 202 507 203 508
rect 203 507 204 508
rect 204 507 205 508
rect 205 507 206 508
rect 206 507 207 508
rect 207 507 208 508
rect 208 507 209 508
rect 226 507 227 508
rect 227 507 228 508
rect 228 507 229 508
rect 229 507 230 508
rect 230 507 231 508
rect 231 507 232 508
rect 232 507 233 508
rect 266 507 267 508
rect 267 507 268 508
rect 268 507 269 508
rect 269 507 270 508
rect 270 507 271 508
rect 271 507 272 508
rect 272 507 273 508
rect 273 507 274 508
rect 274 507 275 508
rect 275 507 276 508
rect 276 507 277 508
rect 277 507 278 508
rect 278 507 279 508
rect 279 507 280 508
rect 280 507 281 508
rect 281 507 282 508
rect 295 507 296 508
rect 296 507 297 508
rect 297 507 298 508
rect 298 507 299 508
rect 299 507 300 508
rect 300 507 301 508
rect 301 507 302 508
rect 302 507 303 508
rect 303 507 304 508
rect 304 507 305 508
rect 305 507 306 508
rect 306 507 307 508
rect 307 507 308 508
rect 308 507 309 508
rect 309 507 310 508
rect 310 507 311 508
rect 311 507 312 508
rect 312 507 313 508
rect 313 507 314 508
rect 314 507 315 508
rect 315 507 316 508
rect 316 507 317 508
rect 317 507 318 508
rect 318 507 319 508
rect 319 507 320 508
rect 320 507 321 508
rect 321 507 322 508
rect 322 507 323 508
rect 323 507 324 508
rect 324 507 325 508
rect 325 507 326 508
rect 326 507 327 508
rect 327 507 328 508
rect 328 507 329 508
rect 329 507 330 508
rect 330 507 331 508
rect 331 507 332 508
rect 332 507 333 508
rect 333 507 334 508
rect 334 507 335 508
rect 335 507 336 508
rect 336 507 337 508
rect 337 507 338 508
rect 338 507 339 508
rect 339 507 340 508
rect 340 507 341 508
rect 341 507 342 508
rect 342 507 343 508
rect 343 507 344 508
rect 344 507 345 508
rect 345 507 346 508
rect 346 507 347 508
rect 347 507 348 508
rect 348 507 349 508
rect 349 507 350 508
rect 350 507 351 508
rect 351 507 352 508
rect 352 507 353 508
rect 353 507 354 508
rect 354 507 355 508
rect 355 507 356 508
rect 356 507 357 508
rect 127 506 128 507
rect 128 506 129 507
rect 129 506 130 507
rect 130 506 131 507
rect 131 506 132 507
rect 132 506 133 507
rect 133 506 134 507
rect 134 506 135 507
rect 135 506 136 507
rect 200 506 201 507
rect 201 506 202 507
rect 202 506 203 507
rect 203 506 204 507
rect 204 506 205 507
rect 205 506 206 507
rect 206 506 207 507
rect 207 506 208 507
rect 208 506 209 507
rect 209 506 210 507
rect 210 506 211 507
rect 227 506 228 507
rect 228 506 229 507
rect 229 506 230 507
rect 230 506 231 507
rect 231 506 232 507
rect 232 506 233 507
rect 233 506 234 507
rect 268 506 269 507
rect 269 506 270 507
rect 270 506 271 507
rect 271 506 272 507
rect 272 506 273 507
rect 273 506 274 507
rect 274 506 275 507
rect 275 506 276 507
rect 276 506 277 507
rect 277 506 278 507
rect 278 506 279 507
rect 279 506 280 507
rect 280 506 281 507
rect 281 506 282 507
rect 282 506 283 507
rect 291 506 292 507
rect 292 506 293 507
rect 293 506 294 507
rect 294 506 295 507
rect 295 506 296 507
rect 296 506 297 507
rect 297 506 298 507
rect 298 506 299 507
rect 299 506 300 507
rect 300 506 301 507
rect 301 506 302 507
rect 302 506 303 507
rect 303 506 304 507
rect 304 506 305 507
rect 305 506 306 507
rect 306 506 307 507
rect 307 506 308 507
rect 308 506 309 507
rect 309 506 310 507
rect 310 506 311 507
rect 311 506 312 507
rect 312 506 313 507
rect 313 506 314 507
rect 314 506 315 507
rect 315 506 316 507
rect 316 506 317 507
rect 317 506 318 507
rect 318 506 319 507
rect 319 506 320 507
rect 320 506 321 507
rect 321 506 322 507
rect 322 506 323 507
rect 323 506 324 507
rect 324 506 325 507
rect 325 506 326 507
rect 326 506 327 507
rect 327 506 328 507
rect 328 506 329 507
rect 329 506 330 507
rect 330 506 331 507
rect 331 506 332 507
rect 332 506 333 507
rect 333 506 334 507
rect 334 506 335 507
rect 335 506 336 507
rect 336 506 337 507
rect 337 506 338 507
rect 338 506 339 507
rect 339 506 340 507
rect 340 506 341 507
rect 341 506 342 507
rect 342 506 343 507
rect 343 506 344 507
rect 344 506 345 507
rect 345 506 346 507
rect 346 506 347 507
rect 347 506 348 507
rect 348 506 349 507
rect 349 506 350 507
rect 350 506 351 507
rect 351 506 352 507
rect 352 506 353 507
rect 353 506 354 507
rect 354 506 355 507
rect 355 506 356 507
rect 356 506 357 507
rect 357 506 358 507
rect 358 506 359 507
rect 359 506 360 507
rect 127 505 128 506
rect 128 505 129 506
rect 129 505 130 506
rect 130 505 131 506
rect 131 505 132 506
rect 132 505 133 506
rect 133 505 134 506
rect 134 505 135 506
rect 135 505 136 506
rect 200 505 201 506
rect 201 505 202 506
rect 202 505 203 506
rect 203 505 204 506
rect 204 505 205 506
rect 205 505 206 506
rect 206 505 207 506
rect 207 505 208 506
rect 208 505 209 506
rect 209 505 210 506
rect 210 505 211 506
rect 211 505 212 506
rect 227 505 228 506
rect 228 505 229 506
rect 229 505 230 506
rect 230 505 231 506
rect 231 505 232 506
rect 232 505 233 506
rect 233 505 234 506
rect 234 505 235 506
rect 269 505 270 506
rect 270 505 271 506
rect 271 505 272 506
rect 272 505 273 506
rect 273 505 274 506
rect 274 505 275 506
rect 275 505 276 506
rect 276 505 277 506
rect 277 505 278 506
rect 278 505 279 506
rect 279 505 280 506
rect 280 505 281 506
rect 281 505 282 506
rect 282 505 283 506
rect 283 505 284 506
rect 284 505 285 506
rect 287 505 288 506
rect 288 505 289 506
rect 289 505 290 506
rect 290 505 291 506
rect 291 505 292 506
rect 292 505 293 506
rect 293 505 294 506
rect 294 505 295 506
rect 295 505 296 506
rect 296 505 297 506
rect 297 505 298 506
rect 298 505 299 506
rect 299 505 300 506
rect 300 505 301 506
rect 301 505 302 506
rect 302 505 303 506
rect 303 505 304 506
rect 304 505 305 506
rect 305 505 306 506
rect 306 505 307 506
rect 307 505 308 506
rect 308 505 309 506
rect 309 505 310 506
rect 310 505 311 506
rect 311 505 312 506
rect 312 505 313 506
rect 313 505 314 506
rect 314 505 315 506
rect 315 505 316 506
rect 316 505 317 506
rect 317 505 318 506
rect 318 505 319 506
rect 319 505 320 506
rect 320 505 321 506
rect 321 505 322 506
rect 322 505 323 506
rect 323 505 324 506
rect 324 505 325 506
rect 325 505 326 506
rect 326 505 327 506
rect 327 505 328 506
rect 328 505 329 506
rect 329 505 330 506
rect 330 505 331 506
rect 331 505 332 506
rect 332 505 333 506
rect 333 505 334 506
rect 334 505 335 506
rect 335 505 336 506
rect 336 505 337 506
rect 337 505 338 506
rect 338 505 339 506
rect 339 505 340 506
rect 340 505 341 506
rect 341 505 342 506
rect 342 505 343 506
rect 343 505 344 506
rect 344 505 345 506
rect 345 505 346 506
rect 346 505 347 506
rect 347 505 348 506
rect 348 505 349 506
rect 349 505 350 506
rect 350 505 351 506
rect 351 505 352 506
rect 352 505 353 506
rect 353 505 354 506
rect 354 505 355 506
rect 355 505 356 506
rect 356 505 357 506
rect 357 505 358 506
rect 358 505 359 506
rect 359 505 360 506
rect 360 505 361 506
rect 361 505 362 506
rect 127 504 128 505
rect 128 504 129 505
rect 129 504 130 505
rect 130 504 131 505
rect 131 504 132 505
rect 132 504 133 505
rect 133 504 134 505
rect 134 504 135 505
rect 135 504 136 505
rect 201 504 202 505
rect 202 504 203 505
rect 203 504 204 505
rect 204 504 205 505
rect 205 504 206 505
rect 206 504 207 505
rect 207 504 208 505
rect 208 504 209 505
rect 209 504 210 505
rect 210 504 211 505
rect 211 504 212 505
rect 212 504 213 505
rect 213 504 214 505
rect 227 504 228 505
rect 228 504 229 505
rect 229 504 230 505
rect 230 504 231 505
rect 231 504 232 505
rect 232 504 233 505
rect 233 504 234 505
rect 234 504 235 505
rect 235 504 236 505
rect 271 504 272 505
rect 272 504 273 505
rect 273 504 274 505
rect 274 504 275 505
rect 275 504 276 505
rect 276 504 277 505
rect 277 504 278 505
rect 278 504 279 505
rect 279 504 280 505
rect 280 504 281 505
rect 281 504 282 505
rect 282 504 283 505
rect 283 504 284 505
rect 284 504 285 505
rect 285 504 286 505
rect 286 504 287 505
rect 287 504 288 505
rect 288 504 289 505
rect 289 504 290 505
rect 290 504 291 505
rect 291 504 292 505
rect 292 504 293 505
rect 293 504 294 505
rect 294 504 295 505
rect 295 504 296 505
rect 296 504 297 505
rect 297 504 298 505
rect 298 504 299 505
rect 299 504 300 505
rect 300 504 301 505
rect 301 504 302 505
rect 302 504 303 505
rect 303 504 304 505
rect 304 504 305 505
rect 305 504 306 505
rect 306 504 307 505
rect 307 504 308 505
rect 308 504 309 505
rect 309 504 310 505
rect 310 504 311 505
rect 311 504 312 505
rect 312 504 313 505
rect 313 504 314 505
rect 314 504 315 505
rect 315 504 316 505
rect 316 504 317 505
rect 317 504 318 505
rect 318 504 319 505
rect 319 504 320 505
rect 320 504 321 505
rect 321 504 322 505
rect 322 504 323 505
rect 323 504 324 505
rect 324 504 325 505
rect 325 504 326 505
rect 326 504 327 505
rect 327 504 328 505
rect 328 504 329 505
rect 329 504 330 505
rect 330 504 331 505
rect 331 504 332 505
rect 332 504 333 505
rect 333 504 334 505
rect 334 504 335 505
rect 335 504 336 505
rect 336 504 337 505
rect 337 504 338 505
rect 338 504 339 505
rect 339 504 340 505
rect 340 504 341 505
rect 341 504 342 505
rect 342 504 343 505
rect 343 504 344 505
rect 344 504 345 505
rect 345 504 346 505
rect 346 504 347 505
rect 347 504 348 505
rect 348 504 349 505
rect 349 504 350 505
rect 350 504 351 505
rect 351 504 352 505
rect 352 504 353 505
rect 353 504 354 505
rect 354 504 355 505
rect 355 504 356 505
rect 356 504 357 505
rect 357 504 358 505
rect 358 504 359 505
rect 359 504 360 505
rect 360 504 361 505
rect 361 504 362 505
rect 362 504 363 505
rect 363 504 364 505
rect 364 504 365 505
rect 127 503 128 504
rect 128 503 129 504
rect 129 503 130 504
rect 130 503 131 504
rect 131 503 132 504
rect 132 503 133 504
rect 133 503 134 504
rect 134 503 135 504
rect 135 503 136 504
rect 201 503 202 504
rect 202 503 203 504
rect 203 503 204 504
rect 204 503 205 504
rect 205 503 206 504
rect 206 503 207 504
rect 207 503 208 504
rect 208 503 209 504
rect 209 503 210 504
rect 210 503 211 504
rect 211 503 212 504
rect 212 503 213 504
rect 213 503 214 504
rect 214 503 215 504
rect 227 503 228 504
rect 228 503 229 504
rect 229 503 230 504
rect 230 503 231 504
rect 231 503 232 504
rect 232 503 233 504
rect 233 503 234 504
rect 234 503 235 504
rect 235 503 236 504
rect 236 503 237 504
rect 273 503 274 504
rect 274 503 275 504
rect 275 503 276 504
rect 276 503 277 504
rect 277 503 278 504
rect 278 503 279 504
rect 279 503 280 504
rect 280 503 281 504
rect 281 503 282 504
rect 282 503 283 504
rect 283 503 284 504
rect 284 503 285 504
rect 285 503 286 504
rect 286 503 287 504
rect 287 503 288 504
rect 288 503 289 504
rect 289 503 290 504
rect 290 503 291 504
rect 291 503 292 504
rect 292 503 293 504
rect 293 503 294 504
rect 294 503 295 504
rect 295 503 296 504
rect 296 503 297 504
rect 297 503 298 504
rect 298 503 299 504
rect 299 503 300 504
rect 300 503 301 504
rect 301 503 302 504
rect 302 503 303 504
rect 303 503 304 504
rect 304 503 305 504
rect 305 503 306 504
rect 306 503 307 504
rect 307 503 308 504
rect 308 503 309 504
rect 309 503 310 504
rect 310 503 311 504
rect 311 503 312 504
rect 312 503 313 504
rect 313 503 314 504
rect 314 503 315 504
rect 315 503 316 504
rect 316 503 317 504
rect 317 503 318 504
rect 318 503 319 504
rect 319 503 320 504
rect 320 503 321 504
rect 321 503 322 504
rect 322 503 323 504
rect 323 503 324 504
rect 324 503 325 504
rect 325 503 326 504
rect 326 503 327 504
rect 327 503 328 504
rect 328 503 329 504
rect 329 503 330 504
rect 330 503 331 504
rect 331 503 332 504
rect 332 503 333 504
rect 333 503 334 504
rect 334 503 335 504
rect 335 503 336 504
rect 336 503 337 504
rect 337 503 338 504
rect 338 503 339 504
rect 339 503 340 504
rect 340 503 341 504
rect 341 503 342 504
rect 342 503 343 504
rect 343 503 344 504
rect 344 503 345 504
rect 345 503 346 504
rect 346 503 347 504
rect 347 503 348 504
rect 348 503 349 504
rect 349 503 350 504
rect 350 503 351 504
rect 351 503 352 504
rect 352 503 353 504
rect 353 503 354 504
rect 354 503 355 504
rect 355 503 356 504
rect 356 503 357 504
rect 357 503 358 504
rect 358 503 359 504
rect 359 503 360 504
rect 360 503 361 504
rect 361 503 362 504
rect 362 503 363 504
rect 363 503 364 504
rect 364 503 365 504
rect 365 503 366 504
rect 366 503 367 504
rect 127 502 128 503
rect 128 502 129 503
rect 129 502 130 503
rect 130 502 131 503
rect 131 502 132 503
rect 132 502 133 503
rect 133 502 134 503
rect 134 502 135 503
rect 135 502 136 503
rect 202 502 203 503
rect 203 502 204 503
rect 204 502 205 503
rect 205 502 206 503
rect 206 502 207 503
rect 207 502 208 503
rect 208 502 209 503
rect 209 502 210 503
rect 210 502 211 503
rect 211 502 212 503
rect 212 502 213 503
rect 213 502 214 503
rect 214 502 215 503
rect 215 502 216 503
rect 216 502 217 503
rect 227 502 228 503
rect 228 502 229 503
rect 229 502 230 503
rect 230 502 231 503
rect 231 502 232 503
rect 232 502 233 503
rect 233 502 234 503
rect 234 502 235 503
rect 235 502 236 503
rect 236 502 237 503
rect 237 502 238 503
rect 274 502 275 503
rect 275 502 276 503
rect 276 502 277 503
rect 277 502 278 503
rect 278 502 279 503
rect 279 502 280 503
rect 280 502 281 503
rect 281 502 282 503
rect 282 502 283 503
rect 283 502 284 503
rect 284 502 285 503
rect 285 502 286 503
rect 286 502 287 503
rect 287 502 288 503
rect 288 502 289 503
rect 289 502 290 503
rect 290 502 291 503
rect 291 502 292 503
rect 292 502 293 503
rect 293 502 294 503
rect 294 502 295 503
rect 295 502 296 503
rect 296 502 297 503
rect 297 502 298 503
rect 298 502 299 503
rect 299 502 300 503
rect 300 502 301 503
rect 301 502 302 503
rect 302 502 303 503
rect 303 502 304 503
rect 304 502 305 503
rect 305 502 306 503
rect 306 502 307 503
rect 307 502 308 503
rect 308 502 309 503
rect 309 502 310 503
rect 310 502 311 503
rect 311 502 312 503
rect 312 502 313 503
rect 313 502 314 503
rect 314 502 315 503
rect 315 502 316 503
rect 316 502 317 503
rect 317 502 318 503
rect 318 502 319 503
rect 319 502 320 503
rect 337 502 338 503
rect 338 502 339 503
rect 339 502 340 503
rect 340 502 341 503
rect 341 502 342 503
rect 342 502 343 503
rect 343 502 344 503
rect 344 502 345 503
rect 345 502 346 503
rect 346 502 347 503
rect 347 502 348 503
rect 348 502 349 503
rect 349 502 350 503
rect 350 502 351 503
rect 351 502 352 503
rect 352 502 353 503
rect 353 502 354 503
rect 354 502 355 503
rect 355 502 356 503
rect 356 502 357 503
rect 357 502 358 503
rect 358 502 359 503
rect 359 502 360 503
rect 360 502 361 503
rect 361 502 362 503
rect 362 502 363 503
rect 363 502 364 503
rect 364 502 365 503
rect 365 502 366 503
rect 366 502 367 503
rect 367 502 368 503
rect 368 502 369 503
rect 128 501 129 502
rect 129 501 130 502
rect 130 501 131 502
rect 131 501 132 502
rect 132 501 133 502
rect 133 501 134 502
rect 134 501 135 502
rect 135 501 136 502
rect 204 501 205 502
rect 205 501 206 502
rect 206 501 207 502
rect 207 501 208 502
rect 208 501 209 502
rect 209 501 210 502
rect 210 501 211 502
rect 211 501 212 502
rect 212 501 213 502
rect 213 501 214 502
rect 214 501 215 502
rect 215 501 216 502
rect 216 501 217 502
rect 217 501 218 502
rect 218 501 219 502
rect 227 501 228 502
rect 228 501 229 502
rect 229 501 230 502
rect 230 501 231 502
rect 231 501 232 502
rect 232 501 233 502
rect 233 501 234 502
rect 234 501 235 502
rect 235 501 236 502
rect 236 501 237 502
rect 237 501 238 502
rect 275 501 276 502
rect 276 501 277 502
rect 277 501 278 502
rect 278 501 279 502
rect 279 501 280 502
rect 280 501 281 502
rect 281 501 282 502
rect 282 501 283 502
rect 283 501 284 502
rect 284 501 285 502
rect 285 501 286 502
rect 286 501 287 502
rect 287 501 288 502
rect 288 501 289 502
rect 289 501 290 502
rect 290 501 291 502
rect 291 501 292 502
rect 292 501 293 502
rect 293 501 294 502
rect 294 501 295 502
rect 295 501 296 502
rect 296 501 297 502
rect 297 501 298 502
rect 298 501 299 502
rect 299 501 300 502
rect 300 501 301 502
rect 301 501 302 502
rect 302 501 303 502
rect 303 501 304 502
rect 304 501 305 502
rect 305 501 306 502
rect 306 501 307 502
rect 307 501 308 502
rect 308 501 309 502
rect 309 501 310 502
rect 310 501 311 502
rect 345 501 346 502
rect 346 501 347 502
rect 347 501 348 502
rect 348 501 349 502
rect 349 501 350 502
rect 350 501 351 502
rect 351 501 352 502
rect 352 501 353 502
rect 353 501 354 502
rect 354 501 355 502
rect 355 501 356 502
rect 356 501 357 502
rect 357 501 358 502
rect 358 501 359 502
rect 359 501 360 502
rect 360 501 361 502
rect 361 501 362 502
rect 362 501 363 502
rect 363 501 364 502
rect 364 501 365 502
rect 365 501 366 502
rect 366 501 367 502
rect 367 501 368 502
rect 368 501 369 502
rect 369 501 370 502
rect 370 501 371 502
rect 128 500 129 501
rect 129 500 130 501
rect 130 500 131 501
rect 131 500 132 501
rect 132 500 133 501
rect 133 500 134 501
rect 134 500 135 501
rect 135 500 136 501
rect 136 500 137 501
rect 206 500 207 501
rect 207 500 208 501
rect 208 500 209 501
rect 209 500 210 501
rect 210 500 211 501
rect 211 500 212 501
rect 212 500 213 501
rect 213 500 214 501
rect 214 500 215 501
rect 215 500 216 501
rect 216 500 217 501
rect 217 500 218 501
rect 218 500 219 501
rect 219 500 220 501
rect 220 500 221 501
rect 226 500 227 501
rect 227 500 228 501
rect 228 500 229 501
rect 229 500 230 501
rect 230 500 231 501
rect 231 500 232 501
rect 232 500 233 501
rect 233 500 234 501
rect 234 500 235 501
rect 235 500 236 501
rect 236 500 237 501
rect 237 500 238 501
rect 238 500 239 501
rect 272 500 273 501
rect 273 500 274 501
rect 274 500 275 501
rect 275 500 276 501
rect 276 500 277 501
rect 277 500 278 501
rect 278 500 279 501
rect 279 500 280 501
rect 280 500 281 501
rect 281 500 282 501
rect 282 500 283 501
rect 283 500 284 501
rect 284 500 285 501
rect 285 500 286 501
rect 286 500 287 501
rect 287 500 288 501
rect 288 500 289 501
rect 289 500 290 501
rect 290 500 291 501
rect 291 500 292 501
rect 292 500 293 501
rect 293 500 294 501
rect 294 500 295 501
rect 295 500 296 501
rect 296 500 297 501
rect 297 500 298 501
rect 298 500 299 501
rect 299 500 300 501
rect 300 500 301 501
rect 301 500 302 501
rect 302 500 303 501
rect 303 500 304 501
rect 304 500 305 501
rect 350 500 351 501
rect 351 500 352 501
rect 352 500 353 501
rect 353 500 354 501
rect 354 500 355 501
rect 355 500 356 501
rect 356 500 357 501
rect 357 500 358 501
rect 358 500 359 501
rect 359 500 360 501
rect 360 500 361 501
rect 361 500 362 501
rect 362 500 363 501
rect 363 500 364 501
rect 364 500 365 501
rect 365 500 366 501
rect 366 500 367 501
rect 367 500 368 501
rect 368 500 369 501
rect 369 500 370 501
rect 370 500 371 501
rect 371 500 372 501
rect 128 499 129 500
rect 129 499 130 500
rect 130 499 131 500
rect 131 499 132 500
rect 132 499 133 500
rect 133 499 134 500
rect 134 499 135 500
rect 135 499 136 500
rect 136 499 137 500
rect 207 499 208 500
rect 208 499 209 500
rect 209 499 210 500
rect 210 499 211 500
rect 211 499 212 500
rect 212 499 213 500
rect 213 499 214 500
rect 214 499 215 500
rect 215 499 216 500
rect 216 499 217 500
rect 217 499 218 500
rect 218 499 219 500
rect 219 499 220 500
rect 220 499 221 500
rect 221 499 222 500
rect 222 499 223 500
rect 223 499 224 500
rect 224 499 225 500
rect 225 499 226 500
rect 226 499 227 500
rect 227 499 228 500
rect 228 499 229 500
rect 229 499 230 500
rect 230 499 231 500
rect 231 499 232 500
rect 232 499 233 500
rect 233 499 234 500
rect 234 499 235 500
rect 235 499 236 500
rect 236 499 237 500
rect 237 499 238 500
rect 238 499 239 500
rect 239 499 240 500
rect 269 499 270 500
rect 270 499 271 500
rect 271 499 272 500
rect 272 499 273 500
rect 273 499 274 500
rect 274 499 275 500
rect 275 499 276 500
rect 276 499 277 500
rect 277 499 278 500
rect 278 499 279 500
rect 279 499 280 500
rect 280 499 281 500
rect 281 499 282 500
rect 282 499 283 500
rect 283 499 284 500
rect 284 499 285 500
rect 285 499 286 500
rect 286 499 287 500
rect 287 499 288 500
rect 288 499 289 500
rect 289 499 290 500
rect 290 499 291 500
rect 291 499 292 500
rect 292 499 293 500
rect 293 499 294 500
rect 294 499 295 500
rect 295 499 296 500
rect 296 499 297 500
rect 297 499 298 500
rect 298 499 299 500
rect 299 499 300 500
rect 354 499 355 500
rect 355 499 356 500
rect 356 499 357 500
rect 357 499 358 500
rect 358 499 359 500
rect 359 499 360 500
rect 360 499 361 500
rect 361 499 362 500
rect 362 499 363 500
rect 363 499 364 500
rect 364 499 365 500
rect 365 499 366 500
rect 366 499 367 500
rect 367 499 368 500
rect 368 499 369 500
rect 369 499 370 500
rect 370 499 371 500
rect 371 499 372 500
rect 372 499 373 500
rect 373 499 374 500
rect 128 498 129 499
rect 129 498 130 499
rect 130 498 131 499
rect 131 498 132 499
rect 132 498 133 499
rect 133 498 134 499
rect 134 498 135 499
rect 135 498 136 499
rect 136 498 137 499
rect 209 498 210 499
rect 210 498 211 499
rect 211 498 212 499
rect 212 498 213 499
rect 213 498 214 499
rect 214 498 215 499
rect 215 498 216 499
rect 216 498 217 499
rect 217 498 218 499
rect 218 498 219 499
rect 219 498 220 499
rect 220 498 221 499
rect 221 498 222 499
rect 222 498 223 499
rect 223 498 224 499
rect 224 498 225 499
rect 225 498 226 499
rect 226 498 227 499
rect 227 498 228 499
rect 228 498 229 499
rect 229 498 230 499
rect 230 498 231 499
rect 231 498 232 499
rect 232 498 233 499
rect 233 498 234 499
rect 234 498 235 499
rect 235 498 236 499
rect 236 498 237 499
rect 237 498 238 499
rect 238 498 239 499
rect 239 498 240 499
rect 267 498 268 499
rect 268 498 269 499
rect 269 498 270 499
rect 270 498 271 499
rect 271 498 272 499
rect 272 498 273 499
rect 273 498 274 499
rect 274 498 275 499
rect 275 498 276 499
rect 276 498 277 499
rect 277 498 278 499
rect 278 498 279 499
rect 279 498 280 499
rect 280 498 281 499
rect 281 498 282 499
rect 282 498 283 499
rect 283 498 284 499
rect 284 498 285 499
rect 285 498 286 499
rect 286 498 287 499
rect 287 498 288 499
rect 288 498 289 499
rect 289 498 290 499
rect 290 498 291 499
rect 291 498 292 499
rect 292 498 293 499
rect 293 498 294 499
rect 294 498 295 499
rect 357 498 358 499
rect 358 498 359 499
rect 359 498 360 499
rect 360 498 361 499
rect 361 498 362 499
rect 362 498 363 499
rect 363 498 364 499
rect 364 498 365 499
rect 365 498 366 499
rect 366 498 367 499
rect 367 498 368 499
rect 368 498 369 499
rect 369 498 370 499
rect 370 498 371 499
rect 371 498 372 499
rect 372 498 373 499
rect 373 498 374 499
rect 374 498 375 499
rect 128 497 129 498
rect 129 497 130 498
rect 130 497 131 498
rect 131 497 132 498
rect 132 497 133 498
rect 133 497 134 498
rect 134 497 135 498
rect 135 497 136 498
rect 136 497 137 498
rect 150 497 151 498
rect 211 497 212 498
rect 212 497 213 498
rect 213 497 214 498
rect 214 497 215 498
rect 215 497 216 498
rect 216 497 217 498
rect 217 497 218 498
rect 218 497 219 498
rect 219 497 220 498
rect 220 497 221 498
rect 221 497 222 498
rect 222 497 223 498
rect 223 497 224 498
rect 224 497 225 498
rect 225 497 226 498
rect 226 497 227 498
rect 227 497 228 498
rect 228 497 229 498
rect 229 497 230 498
rect 230 497 231 498
rect 231 497 232 498
rect 232 497 233 498
rect 233 497 234 498
rect 234 497 235 498
rect 235 497 236 498
rect 236 497 237 498
rect 237 497 238 498
rect 238 497 239 498
rect 239 497 240 498
rect 240 497 241 498
rect 264 497 265 498
rect 265 497 266 498
rect 266 497 267 498
rect 267 497 268 498
rect 268 497 269 498
rect 269 497 270 498
rect 270 497 271 498
rect 271 497 272 498
rect 272 497 273 498
rect 273 497 274 498
rect 274 497 275 498
rect 275 497 276 498
rect 276 497 277 498
rect 277 497 278 498
rect 278 497 279 498
rect 279 497 280 498
rect 280 497 281 498
rect 281 497 282 498
rect 282 497 283 498
rect 283 497 284 498
rect 284 497 285 498
rect 285 497 286 498
rect 286 497 287 498
rect 287 497 288 498
rect 288 497 289 498
rect 289 497 290 498
rect 290 497 291 498
rect 359 497 360 498
rect 360 497 361 498
rect 361 497 362 498
rect 362 497 363 498
rect 363 497 364 498
rect 364 497 365 498
rect 365 497 366 498
rect 366 497 367 498
rect 367 497 368 498
rect 368 497 369 498
rect 369 497 370 498
rect 370 497 371 498
rect 371 497 372 498
rect 372 497 373 498
rect 373 497 374 498
rect 374 497 375 498
rect 375 497 376 498
rect 376 497 377 498
rect 128 496 129 497
rect 129 496 130 497
rect 130 496 131 497
rect 131 496 132 497
rect 132 496 133 497
rect 133 496 134 497
rect 134 496 135 497
rect 135 496 136 497
rect 136 496 137 497
rect 137 496 138 497
rect 151 496 152 497
rect 213 496 214 497
rect 214 496 215 497
rect 215 496 216 497
rect 216 496 217 497
rect 217 496 218 497
rect 218 496 219 497
rect 219 496 220 497
rect 220 496 221 497
rect 221 496 222 497
rect 222 496 223 497
rect 223 496 224 497
rect 224 496 225 497
rect 225 496 226 497
rect 226 496 227 497
rect 227 496 228 497
rect 228 496 229 497
rect 229 496 230 497
rect 230 496 231 497
rect 231 496 232 497
rect 232 496 233 497
rect 233 496 234 497
rect 234 496 235 497
rect 235 496 236 497
rect 236 496 237 497
rect 237 496 238 497
rect 238 496 239 497
rect 239 496 240 497
rect 240 496 241 497
rect 262 496 263 497
rect 263 496 264 497
rect 264 496 265 497
rect 265 496 266 497
rect 266 496 267 497
rect 267 496 268 497
rect 268 496 269 497
rect 269 496 270 497
rect 270 496 271 497
rect 271 496 272 497
rect 272 496 273 497
rect 273 496 274 497
rect 274 496 275 497
rect 275 496 276 497
rect 276 496 277 497
rect 277 496 278 497
rect 278 496 279 497
rect 279 496 280 497
rect 280 496 281 497
rect 281 496 282 497
rect 282 496 283 497
rect 283 496 284 497
rect 284 496 285 497
rect 285 496 286 497
rect 286 496 287 497
rect 287 496 288 497
rect 362 496 363 497
rect 363 496 364 497
rect 364 496 365 497
rect 365 496 366 497
rect 366 496 367 497
rect 367 496 368 497
rect 368 496 369 497
rect 369 496 370 497
rect 370 496 371 497
rect 371 496 372 497
rect 372 496 373 497
rect 373 496 374 497
rect 374 496 375 497
rect 375 496 376 497
rect 376 496 377 497
rect 377 496 378 497
rect 378 496 379 497
rect 129 495 130 496
rect 130 495 131 496
rect 131 495 132 496
rect 132 495 133 496
rect 133 495 134 496
rect 134 495 135 496
rect 135 495 136 496
rect 136 495 137 496
rect 137 495 138 496
rect 151 495 152 496
rect 152 495 153 496
rect 215 495 216 496
rect 216 495 217 496
rect 217 495 218 496
rect 218 495 219 496
rect 219 495 220 496
rect 220 495 221 496
rect 221 495 222 496
rect 222 495 223 496
rect 223 495 224 496
rect 224 495 225 496
rect 225 495 226 496
rect 226 495 227 496
rect 227 495 228 496
rect 228 495 229 496
rect 229 495 230 496
rect 230 495 231 496
rect 231 495 232 496
rect 232 495 233 496
rect 233 495 234 496
rect 234 495 235 496
rect 235 495 236 496
rect 236 495 237 496
rect 237 495 238 496
rect 238 495 239 496
rect 239 495 240 496
rect 240 495 241 496
rect 259 495 260 496
rect 260 495 261 496
rect 261 495 262 496
rect 262 495 263 496
rect 263 495 264 496
rect 264 495 265 496
rect 265 495 266 496
rect 266 495 267 496
rect 267 495 268 496
rect 268 495 269 496
rect 269 495 270 496
rect 270 495 271 496
rect 271 495 272 496
rect 272 495 273 496
rect 273 495 274 496
rect 274 495 275 496
rect 275 495 276 496
rect 276 495 277 496
rect 277 495 278 496
rect 278 495 279 496
rect 279 495 280 496
rect 280 495 281 496
rect 281 495 282 496
rect 282 495 283 496
rect 283 495 284 496
rect 364 495 365 496
rect 365 495 366 496
rect 366 495 367 496
rect 367 495 368 496
rect 368 495 369 496
rect 369 495 370 496
rect 370 495 371 496
rect 371 495 372 496
rect 372 495 373 496
rect 373 495 374 496
rect 374 495 375 496
rect 375 495 376 496
rect 376 495 377 496
rect 377 495 378 496
rect 378 495 379 496
rect 379 495 380 496
rect 129 494 130 495
rect 130 494 131 495
rect 131 494 132 495
rect 132 494 133 495
rect 133 494 134 495
rect 134 494 135 495
rect 135 494 136 495
rect 136 494 137 495
rect 137 494 138 495
rect 151 494 152 495
rect 152 494 153 495
rect 217 494 218 495
rect 218 494 219 495
rect 219 494 220 495
rect 220 494 221 495
rect 221 494 222 495
rect 222 494 223 495
rect 223 494 224 495
rect 224 494 225 495
rect 225 494 226 495
rect 226 494 227 495
rect 227 494 228 495
rect 228 494 229 495
rect 229 494 230 495
rect 230 494 231 495
rect 231 494 232 495
rect 232 494 233 495
rect 233 494 234 495
rect 234 494 235 495
rect 235 494 236 495
rect 236 494 237 495
rect 237 494 238 495
rect 238 494 239 495
rect 239 494 240 495
rect 240 494 241 495
rect 257 494 258 495
rect 258 494 259 495
rect 259 494 260 495
rect 260 494 261 495
rect 261 494 262 495
rect 262 494 263 495
rect 263 494 264 495
rect 264 494 265 495
rect 265 494 266 495
rect 266 494 267 495
rect 267 494 268 495
rect 268 494 269 495
rect 269 494 270 495
rect 270 494 271 495
rect 271 494 272 495
rect 272 494 273 495
rect 273 494 274 495
rect 274 494 275 495
rect 275 494 276 495
rect 276 494 277 495
rect 277 494 278 495
rect 278 494 279 495
rect 279 494 280 495
rect 280 494 281 495
rect 366 494 367 495
rect 367 494 368 495
rect 368 494 369 495
rect 369 494 370 495
rect 370 494 371 495
rect 371 494 372 495
rect 372 494 373 495
rect 373 494 374 495
rect 374 494 375 495
rect 375 494 376 495
rect 376 494 377 495
rect 377 494 378 495
rect 378 494 379 495
rect 379 494 380 495
rect 380 494 381 495
rect 381 494 382 495
rect 129 493 130 494
rect 130 493 131 494
rect 131 493 132 494
rect 132 493 133 494
rect 133 493 134 494
rect 134 493 135 494
rect 135 493 136 494
rect 136 493 137 494
rect 137 493 138 494
rect 152 493 153 494
rect 153 493 154 494
rect 219 493 220 494
rect 220 493 221 494
rect 221 493 222 494
rect 222 493 223 494
rect 223 493 224 494
rect 224 493 225 494
rect 225 493 226 494
rect 226 493 227 494
rect 227 493 228 494
rect 228 493 229 494
rect 229 493 230 494
rect 230 493 231 494
rect 231 493 232 494
rect 232 493 233 494
rect 233 493 234 494
rect 234 493 235 494
rect 235 493 236 494
rect 236 493 237 494
rect 237 493 238 494
rect 238 493 239 494
rect 239 493 240 494
rect 240 493 241 494
rect 254 493 255 494
rect 255 493 256 494
rect 256 493 257 494
rect 257 493 258 494
rect 258 493 259 494
rect 259 493 260 494
rect 260 493 261 494
rect 261 493 262 494
rect 262 493 263 494
rect 263 493 264 494
rect 264 493 265 494
rect 265 493 266 494
rect 266 493 267 494
rect 267 493 268 494
rect 268 493 269 494
rect 269 493 270 494
rect 270 493 271 494
rect 271 493 272 494
rect 272 493 273 494
rect 273 493 274 494
rect 274 493 275 494
rect 275 493 276 494
rect 276 493 277 494
rect 277 493 278 494
rect 368 493 369 494
rect 369 493 370 494
rect 370 493 371 494
rect 371 493 372 494
rect 372 493 373 494
rect 373 493 374 494
rect 374 493 375 494
rect 375 493 376 494
rect 376 493 377 494
rect 377 493 378 494
rect 378 493 379 494
rect 379 493 380 494
rect 380 493 381 494
rect 381 493 382 494
rect 382 493 383 494
rect 130 492 131 493
rect 131 492 132 493
rect 132 492 133 493
rect 133 492 134 493
rect 134 492 135 493
rect 135 492 136 493
rect 136 492 137 493
rect 137 492 138 493
rect 138 492 139 493
rect 152 492 153 493
rect 153 492 154 493
rect 222 492 223 493
rect 223 492 224 493
rect 224 492 225 493
rect 225 492 226 493
rect 226 492 227 493
rect 227 492 228 493
rect 228 492 229 493
rect 229 492 230 493
rect 230 492 231 493
rect 231 492 232 493
rect 232 492 233 493
rect 233 492 234 493
rect 234 492 235 493
rect 235 492 236 493
rect 236 492 237 493
rect 237 492 238 493
rect 238 492 239 493
rect 239 492 240 493
rect 240 492 241 493
rect 252 492 253 493
rect 253 492 254 493
rect 254 492 255 493
rect 255 492 256 493
rect 256 492 257 493
rect 257 492 258 493
rect 258 492 259 493
rect 259 492 260 493
rect 260 492 261 493
rect 261 492 262 493
rect 262 492 263 493
rect 263 492 264 493
rect 264 492 265 493
rect 265 492 266 493
rect 266 492 267 493
rect 267 492 268 493
rect 268 492 269 493
rect 269 492 270 493
rect 270 492 271 493
rect 271 492 272 493
rect 272 492 273 493
rect 273 492 274 493
rect 274 492 275 493
rect 369 492 370 493
rect 370 492 371 493
rect 371 492 372 493
rect 372 492 373 493
rect 373 492 374 493
rect 374 492 375 493
rect 375 492 376 493
rect 376 492 377 493
rect 377 492 378 493
rect 378 492 379 493
rect 379 492 380 493
rect 380 492 381 493
rect 381 492 382 493
rect 382 492 383 493
rect 383 492 384 493
rect 384 492 385 493
rect 130 491 131 492
rect 131 491 132 492
rect 132 491 133 492
rect 133 491 134 492
rect 134 491 135 492
rect 135 491 136 492
rect 136 491 137 492
rect 137 491 138 492
rect 138 491 139 492
rect 152 491 153 492
rect 153 491 154 492
rect 154 491 155 492
rect 224 491 225 492
rect 225 491 226 492
rect 226 491 227 492
rect 227 491 228 492
rect 228 491 229 492
rect 229 491 230 492
rect 230 491 231 492
rect 231 491 232 492
rect 232 491 233 492
rect 233 491 234 492
rect 234 491 235 492
rect 235 491 236 492
rect 236 491 237 492
rect 237 491 238 492
rect 238 491 239 492
rect 239 491 240 492
rect 250 491 251 492
rect 251 491 252 492
rect 252 491 253 492
rect 253 491 254 492
rect 254 491 255 492
rect 255 491 256 492
rect 256 491 257 492
rect 257 491 258 492
rect 258 491 259 492
rect 259 491 260 492
rect 260 491 261 492
rect 261 491 262 492
rect 262 491 263 492
rect 263 491 264 492
rect 264 491 265 492
rect 265 491 266 492
rect 266 491 267 492
rect 267 491 268 492
rect 268 491 269 492
rect 269 491 270 492
rect 270 491 271 492
rect 271 491 272 492
rect 371 491 372 492
rect 372 491 373 492
rect 373 491 374 492
rect 374 491 375 492
rect 375 491 376 492
rect 376 491 377 492
rect 377 491 378 492
rect 378 491 379 492
rect 379 491 380 492
rect 380 491 381 492
rect 381 491 382 492
rect 382 491 383 492
rect 383 491 384 492
rect 384 491 385 492
rect 385 491 386 492
rect 386 491 387 492
rect 130 490 131 491
rect 131 490 132 491
rect 132 490 133 491
rect 133 490 134 491
rect 134 490 135 491
rect 135 490 136 491
rect 136 490 137 491
rect 137 490 138 491
rect 138 490 139 491
rect 139 490 140 491
rect 153 490 154 491
rect 154 490 155 491
rect 227 490 228 491
rect 228 490 229 491
rect 229 490 230 491
rect 230 490 231 491
rect 231 490 232 491
rect 232 490 233 491
rect 233 490 234 491
rect 234 490 235 491
rect 235 490 236 491
rect 236 490 237 491
rect 237 490 238 491
rect 238 490 239 491
rect 248 490 249 491
rect 249 490 250 491
rect 250 490 251 491
rect 251 490 252 491
rect 252 490 253 491
rect 253 490 254 491
rect 254 490 255 491
rect 255 490 256 491
rect 256 490 257 491
rect 257 490 258 491
rect 258 490 259 491
rect 259 490 260 491
rect 260 490 261 491
rect 261 490 262 491
rect 262 490 263 491
rect 263 490 264 491
rect 264 490 265 491
rect 265 490 266 491
rect 266 490 267 491
rect 267 490 268 491
rect 268 490 269 491
rect 372 490 373 491
rect 373 490 374 491
rect 374 490 375 491
rect 375 490 376 491
rect 376 490 377 491
rect 377 490 378 491
rect 378 490 379 491
rect 379 490 380 491
rect 380 490 381 491
rect 381 490 382 491
rect 382 490 383 491
rect 383 490 384 491
rect 384 490 385 491
rect 385 490 386 491
rect 386 490 387 491
rect 387 490 388 491
rect 131 489 132 490
rect 132 489 133 490
rect 133 489 134 490
rect 134 489 135 490
rect 135 489 136 490
rect 136 489 137 490
rect 137 489 138 490
rect 138 489 139 490
rect 139 489 140 490
rect 153 489 154 490
rect 154 489 155 490
rect 155 489 156 490
rect 234 489 235 490
rect 246 489 247 490
rect 247 489 248 490
rect 248 489 249 490
rect 249 489 250 490
rect 250 489 251 490
rect 251 489 252 490
rect 252 489 253 490
rect 253 489 254 490
rect 254 489 255 490
rect 255 489 256 490
rect 256 489 257 490
rect 257 489 258 490
rect 258 489 259 490
rect 259 489 260 490
rect 260 489 261 490
rect 261 489 262 490
rect 262 489 263 490
rect 263 489 264 490
rect 264 489 265 490
rect 265 489 266 490
rect 266 489 267 490
rect 374 489 375 490
rect 375 489 376 490
rect 376 489 377 490
rect 377 489 378 490
rect 378 489 379 490
rect 379 489 380 490
rect 380 489 381 490
rect 381 489 382 490
rect 382 489 383 490
rect 383 489 384 490
rect 384 489 385 490
rect 385 489 386 490
rect 386 489 387 490
rect 387 489 388 490
rect 388 489 389 490
rect 389 489 390 490
rect 131 488 132 489
rect 132 488 133 489
rect 133 488 134 489
rect 134 488 135 489
rect 135 488 136 489
rect 136 488 137 489
rect 137 488 138 489
rect 138 488 139 489
rect 139 488 140 489
rect 153 488 154 489
rect 154 488 155 489
rect 155 488 156 489
rect 156 488 157 489
rect 243 488 244 489
rect 244 488 245 489
rect 245 488 246 489
rect 246 488 247 489
rect 247 488 248 489
rect 248 488 249 489
rect 249 488 250 489
rect 250 488 251 489
rect 251 488 252 489
rect 252 488 253 489
rect 253 488 254 489
rect 254 488 255 489
rect 255 488 256 489
rect 256 488 257 489
rect 257 488 258 489
rect 258 488 259 489
rect 259 488 260 489
rect 260 488 261 489
rect 261 488 262 489
rect 262 488 263 489
rect 263 488 264 489
rect 376 488 377 489
rect 377 488 378 489
rect 378 488 379 489
rect 379 488 380 489
rect 380 488 381 489
rect 381 488 382 489
rect 382 488 383 489
rect 383 488 384 489
rect 384 488 385 489
rect 385 488 386 489
rect 386 488 387 489
rect 387 488 388 489
rect 388 488 389 489
rect 389 488 390 489
rect 390 488 391 489
rect 131 487 132 488
rect 132 487 133 488
rect 133 487 134 488
rect 134 487 135 488
rect 135 487 136 488
rect 136 487 137 488
rect 137 487 138 488
rect 138 487 139 488
rect 139 487 140 488
rect 140 487 141 488
rect 154 487 155 488
rect 155 487 156 488
rect 156 487 157 488
rect 241 487 242 488
rect 242 487 243 488
rect 243 487 244 488
rect 244 487 245 488
rect 245 487 246 488
rect 246 487 247 488
rect 247 487 248 488
rect 248 487 249 488
rect 249 487 250 488
rect 250 487 251 488
rect 251 487 252 488
rect 252 487 253 488
rect 253 487 254 488
rect 254 487 255 488
rect 255 487 256 488
rect 256 487 257 488
rect 257 487 258 488
rect 258 487 259 488
rect 259 487 260 488
rect 260 487 261 488
rect 261 487 262 488
rect 377 487 378 488
rect 378 487 379 488
rect 379 487 380 488
rect 380 487 381 488
rect 381 487 382 488
rect 382 487 383 488
rect 383 487 384 488
rect 384 487 385 488
rect 385 487 386 488
rect 386 487 387 488
rect 387 487 388 488
rect 388 487 389 488
rect 389 487 390 488
rect 390 487 391 488
rect 391 487 392 488
rect 392 487 393 488
rect 132 486 133 487
rect 133 486 134 487
rect 134 486 135 487
rect 135 486 136 487
rect 136 486 137 487
rect 137 486 138 487
rect 138 486 139 487
rect 139 486 140 487
rect 140 486 141 487
rect 154 486 155 487
rect 155 486 156 487
rect 156 486 157 487
rect 157 486 158 487
rect 240 486 241 487
rect 241 486 242 487
rect 242 486 243 487
rect 243 486 244 487
rect 244 486 245 487
rect 245 486 246 487
rect 246 486 247 487
rect 247 486 248 487
rect 248 486 249 487
rect 249 486 250 487
rect 250 486 251 487
rect 251 486 252 487
rect 252 486 253 487
rect 253 486 254 487
rect 254 486 255 487
rect 255 486 256 487
rect 256 486 257 487
rect 257 486 258 487
rect 258 486 259 487
rect 379 486 380 487
rect 380 486 381 487
rect 381 486 382 487
rect 382 486 383 487
rect 383 486 384 487
rect 384 486 385 487
rect 385 486 386 487
rect 386 486 387 487
rect 387 486 388 487
rect 388 486 389 487
rect 389 486 390 487
rect 390 486 391 487
rect 391 486 392 487
rect 392 486 393 487
rect 393 486 394 487
rect 132 485 133 486
rect 133 485 134 486
rect 134 485 135 486
rect 135 485 136 486
rect 136 485 137 486
rect 137 485 138 486
rect 138 485 139 486
rect 139 485 140 486
rect 140 485 141 486
rect 141 485 142 486
rect 154 485 155 486
rect 155 485 156 486
rect 156 485 157 486
rect 157 485 158 486
rect 238 485 239 486
rect 239 485 240 486
rect 240 485 241 486
rect 241 485 242 486
rect 242 485 243 486
rect 243 485 244 486
rect 244 485 245 486
rect 245 485 246 486
rect 246 485 247 486
rect 247 485 248 486
rect 248 485 249 486
rect 249 485 250 486
rect 250 485 251 486
rect 251 485 252 486
rect 252 485 253 486
rect 253 485 254 486
rect 254 485 255 486
rect 255 485 256 486
rect 256 485 257 486
rect 380 485 381 486
rect 381 485 382 486
rect 382 485 383 486
rect 383 485 384 486
rect 384 485 385 486
rect 385 485 386 486
rect 386 485 387 486
rect 387 485 388 486
rect 388 485 389 486
rect 389 485 390 486
rect 390 485 391 486
rect 391 485 392 486
rect 392 485 393 486
rect 393 485 394 486
rect 394 485 395 486
rect 395 485 396 486
rect 133 484 134 485
rect 134 484 135 485
rect 135 484 136 485
rect 136 484 137 485
rect 137 484 138 485
rect 138 484 139 485
rect 139 484 140 485
rect 140 484 141 485
rect 141 484 142 485
rect 155 484 156 485
rect 156 484 157 485
rect 157 484 158 485
rect 158 484 159 485
rect 236 484 237 485
rect 237 484 238 485
rect 238 484 239 485
rect 239 484 240 485
rect 240 484 241 485
rect 241 484 242 485
rect 242 484 243 485
rect 243 484 244 485
rect 244 484 245 485
rect 245 484 246 485
rect 246 484 247 485
rect 247 484 248 485
rect 248 484 249 485
rect 249 484 250 485
rect 250 484 251 485
rect 251 484 252 485
rect 252 484 253 485
rect 253 484 254 485
rect 254 484 255 485
rect 382 484 383 485
rect 383 484 384 485
rect 384 484 385 485
rect 385 484 386 485
rect 386 484 387 485
rect 387 484 388 485
rect 388 484 389 485
rect 389 484 390 485
rect 390 484 391 485
rect 391 484 392 485
rect 392 484 393 485
rect 393 484 394 485
rect 394 484 395 485
rect 395 484 396 485
rect 396 484 397 485
rect 133 483 134 484
rect 134 483 135 484
rect 135 483 136 484
rect 136 483 137 484
rect 137 483 138 484
rect 138 483 139 484
rect 139 483 140 484
rect 140 483 141 484
rect 141 483 142 484
rect 155 483 156 484
rect 156 483 157 484
rect 157 483 158 484
rect 158 483 159 484
rect 234 483 235 484
rect 235 483 236 484
rect 236 483 237 484
rect 237 483 238 484
rect 238 483 239 484
rect 239 483 240 484
rect 240 483 241 484
rect 241 483 242 484
rect 242 483 243 484
rect 243 483 244 484
rect 244 483 245 484
rect 245 483 246 484
rect 246 483 247 484
rect 247 483 248 484
rect 248 483 249 484
rect 249 483 250 484
rect 250 483 251 484
rect 251 483 252 484
rect 252 483 253 484
rect 384 483 385 484
rect 385 483 386 484
rect 386 483 387 484
rect 387 483 388 484
rect 388 483 389 484
rect 389 483 390 484
rect 390 483 391 484
rect 391 483 392 484
rect 392 483 393 484
rect 393 483 394 484
rect 394 483 395 484
rect 395 483 396 484
rect 396 483 397 484
rect 397 483 398 484
rect 398 483 399 484
rect 133 482 134 483
rect 134 482 135 483
rect 135 482 136 483
rect 136 482 137 483
rect 137 482 138 483
rect 138 482 139 483
rect 139 482 140 483
rect 140 482 141 483
rect 141 482 142 483
rect 142 482 143 483
rect 155 482 156 483
rect 156 482 157 483
rect 157 482 158 483
rect 158 482 159 483
rect 159 482 160 483
rect 232 482 233 483
rect 233 482 234 483
rect 234 482 235 483
rect 235 482 236 483
rect 236 482 237 483
rect 237 482 238 483
rect 238 482 239 483
rect 239 482 240 483
rect 240 482 241 483
rect 241 482 242 483
rect 242 482 243 483
rect 243 482 244 483
rect 244 482 245 483
rect 245 482 246 483
rect 246 482 247 483
rect 247 482 248 483
rect 248 482 249 483
rect 249 482 250 483
rect 385 482 386 483
rect 386 482 387 483
rect 387 482 388 483
rect 388 482 389 483
rect 389 482 390 483
rect 390 482 391 483
rect 391 482 392 483
rect 392 482 393 483
rect 393 482 394 483
rect 394 482 395 483
rect 395 482 396 483
rect 396 482 397 483
rect 397 482 398 483
rect 398 482 399 483
rect 399 482 400 483
rect 134 481 135 482
rect 135 481 136 482
rect 136 481 137 482
rect 137 481 138 482
rect 138 481 139 482
rect 139 481 140 482
rect 140 481 141 482
rect 141 481 142 482
rect 142 481 143 482
rect 156 481 157 482
rect 157 481 158 482
rect 158 481 159 482
rect 159 481 160 482
rect 230 481 231 482
rect 231 481 232 482
rect 232 481 233 482
rect 233 481 234 482
rect 234 481 235 482
rect 235 481 236 482
rect 236 481 237 482
rect 237 481 238 482
rect 238 481 239 482
rect 239 481 240 482
rect 240 481 241 482
rect 241 481 242 482
rect 242 481 243 482
rect 243 481 244 482
rect 244 481 245 482
rect 245 481 246 482
rect 246 481 247 482
rect 247 481 248 482
rect 387 481 388 482
rect 388 481 389 482
rect 389 481 390 482
rect 390 481 391 482
rect 391 481 392 482
rect 392 481 393 482
rect 393 481 394 482
rect 394 481 395 482
rect 395 481 396 482
rect 396 481 397 482
rect 397 481 398 482
rect 398 481 399 482
rect 399 481 400 482
rect 400 481 401 482
rect 401 481 402 482
rect 134 480 135 481
rect 135 480 136 481
rect 136 480 137 481
rect 137 480 138 481
rect 138 480 139 481
rect 139 480 140 481
rect 140 480 141 481
rect 141 480 142 481
rect 142 480 143 481
rect 156 480 157 481
rect 157 480 158 481
rect 158 480 159 481
rect 159 480 160 481
rect 160 480 161 481
rect 228 480 229 481
rect 229 480 230 481
rect 230 480 231 481
rect 231 480 232 481
rect 232 480 233 481
rect 233 480 234 481
rect 234 480 235 481
rect 235 480 236 481
rect 236 480 237 481
rect 237 480 238 481
rect 238 480 239 481
rect 239 480 240 481
rect 240 480 241 481
rect 241 480 242 481
rect 242 480 243 481
rect 243 480 244 481
rect 244 480 245 481
rect 245 480 246 481
rect 388 480 389 481
rect 389 480 390 481
rect 390 480 391 481
rect 391 480 392 481
rect 392 480 393 481
rect 393 480 394 481
rect 394 480 395 481
rect 395 480 396 481
rect 396 480 397 481
rect 397 480 398 481
rect 398 480 399 481
rect 399 480 400 481
rect 400 480 401 481
rect 401 480 402 481
rect 402 480 403 481
rect 134 479 135 480
rect 135 479 136 480
rect 136 479 137 480
rect 137 479 138 480
rect 138 479 139 480
rect 139 479 140 480
rect 140 479 141 480
rect 141 479 142 480
rect 142 479 143 480
rect 143 479 144 480
rect 156 479 157 480
rect 157 479 158 480
rect 158 479 159 480
rect 159 479 160 480
rect 160 479 161 480
rect 226 479 227 480
rect 227 479 228 480
rect 228 479 229 480
rect 229 479 230 480
rect 230 479 231 480
rect 231 479 232 480
rect 232 479 233 480
rect 233 479 234 480
rect 234 479 235 480
rect 235 479 236 480
rect 236 479 237 480
rect 237 479 238 480
rect 238 479 239 480
rect 239 479 240 480
rect 240 479 241 480
rect 241 479 242 480
rect 242 479 243 480
rect 243 479 244 480
rect 390 479 391 480
rect 391 479 392 480
rect 392 479 393 480
rect 393 479 394 480
rect 394 479 395 480
rect 395 479 396 480
rect 396 479 397 480
rect 397 479 398 480
rect 398 479 399 480
rect 399 479 400 480
rect 400 479 401 480
rect 401 479 402 480
rect 402 479 403 480
rect 403 479 404 480
rect 404 479 405 480
rect 135 478 136 479
rect 136 478 137 479
rect 137 478 138 479
rect 138 478 139 479
rect 139 478 140 479
rect 140 478 141 479
rect 141 478 142 479
rect 142 478 143 479
rect 143 478 144 479
rect 157 478 158 479
rect 158 478 159 479
rect 159 478 160 479
rect 160 478 161 479
rect 161 478 162 479
rect 225 478 226 479
rect 226 478 227 479
rect 227 478 228 479
rect 228 478 229 479
rect 229 478 230 479
rect 230 478 231 479
rect 231 478 232 479
rect 232 478 233 479
rect 233 478 234 479
rect 234 478 235 479
rect 235 478 236 479
rect 236 478 237 479
rect 237 478 238 479
rect 238 478 239 479
rect 239 478 240 479
rect 240 478 241 479
rect 241 478 242 479
rect 391 478 392 479
rect 392 478 393 479
rect 393 478 394 479
rect 394 478 395 479
rect 395 478 396 479
rect 396 478 397 479
rect 397 478 398 479
rect 398 478 399 479
rect 399 478 400 479
rect 400 478 401 479
rect 401 478 402 479
rect 402 478 403 479
rect 403 478 404 479
rect 404 478 405 479
rect 405 478 406 479
rect 135 477 136 478
rect 136 477 137 478
rect 137 477 138 478
rect 138 477 139 478
rect 139 477 140 478
rect 140 477 141 478
rect 141 477 142 478
rect 142 477 143 478
rect 143 477 144 478
rect 157 477 158 478
rect 158 477 159 478
rect 159 477 160 478
rect 160 477 161 478
rect 161 477 162 478
rect 223 477 224 478
rect 224 477 225 478
rect 225 477 226 478
rect 226 477 227 478
rect 227 477 228 478
rect 228 477 229 478
rect 229 477 230 478
rect 230 477 231 478
rect 231 477 232 478
rect 232 477 233 478
rect 233 477 234 478
rect 234 477 235 478
rect 235 477 236 478
rect 236 477 237 478
rect 237 477 238 478
rect 238 477 239 478
rect 239 477 240 478
rect 393 477 394 478
rect 394 477 395 478
rect 395 477 396 478
rect 396 477 397 478
rect 397 477 398 478
rect 398 477 399 478
rect 399 477 400 478
rect 400 477 401 478
rect 401 477 402 478
rect 402 477 403 478
rect 403 477 404 478
rect 404 477 405 478
rect 405 477 406 478
rect 406 477 407 478
rect 407 477 408 478
rect 135 476 136 477
rect 136 476 137 477
rect 137 476 138 477
rect 138 476 139 477
rect 139 476 140 477
rect 140 476 141 477
rect 141 476 142 477
rect 142 476 143 477
rect 143 476 144 477
rect 144 476 145 477
rect 157 476 158 477
rect 158 476 159 477
rect 159 476 160 477
rect 160 476 161 477
rect 161 476 162 477
rect 221 476 222 477
rect 222 476 223 477
rect 223 476 224 477
rect 224 476 225 477
rect 225 476 226 477
rect 226 476 227 477
rect 227 476 228 477
rect 228 476 229 477
rect 229 476 230 477
rect 230 476 231 477
rect 231 476 232 477
rect 232 476 233 477
rect 233 476 234 477
rect 234 476 235 477
rect 235 476 236 477
rect 236 476 237 477
rect 237 476 238 477
rect 394 476 395 477
rect 395 476 396 477
rect 396 476 397 477
rect 397 476 398 477
rect 398 476 399 477
rect 399 476 400 477
rect 400 476 401 477
rect 401 476 402 477
rect 402 476 403 477
rect 403 476 404 477
rect 404 476 405 477
rect 405 476 406 477
rect 406 476 407 477
rect 407 476 408 477
rect 408 476 409 477
rect 136 475 137 476
rect 137 475 138 476
rect 138 475 139 476
rect 139 475 140 476
rect 140 475 141 476
rect 141 475 142 476
rect 142 475 143 476
rect 143 475 144 476
rect 144 475 145 476
rect 158 475 159 476
rect 159 475 160 476
rect 160 475 161 476
rect 161 475 162 476
rect 162 475 163 476
rect 219 475 220 476
rect 220 475 221 476
rect 221 475 222 476
rect 222 475 223 476
rect 223 475 224 476
rect 224 475 225 476
rect 225 475 226 476
rect 226 475 227 476
rect 227 475 228 476
rect 228 475 229 476
rect 229 475 230 476
rect 230 475 231 476
rect 231 475 232 476
rect 232 475 233 476
rect 233 475 234 476
rect 234 475 235 476
rect 235 475 236 476
rect 396 475 397 476
rect 397 475 398 476
rect 398 475 399 476
rect 399 475 400 476
rect 400 475 401 476
rect 401 475 402 476
rect 402 475 403 476
rect 403 475 404 476
rect 404 475 405 476
rect 405 475 406 476
rect 406 475 407 476
rect 407 475 408 476
rect 408 475 409 476
rect 409 475 410 476
rect 136 474 137 475
rect 137 474 138 475
rect 138 474 139 475
rect 139 474 140 475
rect 140 474 141 475
rect 141 474 142 475
rect 142 474 143 475
rect 143 474 144 475
rect 144 474 145 475
rect 158 474 159 475
rect 159 474 160 475
rect 160 474 161 475
rect 161 474 162 475
rect 162 474 163 475
rect 218 474 219 475
rect 219 474 220 475
rect 220 474 221 475
rect 221 474 222 475
rect 222 474 223 475
rect 223 474 224 475
rect 224 474 225 475
rect 225 474 226 475
rect 226 474 227 475
rect 227 474 228 475
rect 228 474 229 475
rect 229 474 230 475
rect 230 474 231 475
rect 231 474 232 475
rect 232 474 233 475
rect 233 474 234 475
rect 234 474 235 475
rect 397 474 398 475
rect 398 474 399 475
rect 399 474 400 475
rect 400 474 401 475
rect 401 474 402 475
rect 402 474 403 475
rect 403 474 404 475
rect 404 474 405 475
rect 405 474 406 475
rect 406 474 407 475
rect 407 474 408 475
rect 408 474 409 475
rect 409 474 410 475
rect 410 474 411 475
rect 411 474 412 475
rect 136 473 137 474
rect 137 473 138 474
rect 138 473 139 474
rect 139 473 140 474
rect 140 473 141 474
rect 141 473 142 474
rect 142 473 143 474
rect 143 473 144 474
rect 144 473 145 474
rect 145 473 146 474
rect 158 473 159 474
rect 159 473 160 474
rect 160 473 161 474
rect 161 473 162 474
rect 162 473 163 474
rect 163 473 164 474
rect 216 473 217 474
rect 217 473 218 474
rect 218 473 219 474
rect 219 473 220 474
rect 220 473 221 474
rect 221 473 222 474
rect 222 473 223 474
rect 223 473 224 474
rect 224 473 225 474
rect 225 473 226 474
rect 226 473 227 474
rect 227 473 228 474
rect 228 473 229 474
rect 229 473 230 474
rect 230 473 231 474
rect 231 473 232 474
rect 232 473 233 474
rect 399 473 400 474
rect 400 473 401 474
rect 401 473 402 474
rect 402 473 403 474
rect 403 473 404 474
rect 404 473 405 474
rect 405 473 406 474
rect 406 473 407 474
rect 407 473 408 474
rect 408 473 409 474
rect 409 473 410 474
rect 410 473 411 474
rect 411 473 412 474
rect 412 473 413 474
rect 137 472 138 473
rect 138 472 139 473
rect 139 472 140 473
rect 140 472 141 473
rect 141 472 142 473
rect 142 472 143 473
rect 143 472 144 473
rect 144 472 145 473
rect 145 472 146 473
rect 159 472 160 473
rect 160 472 161 473
rect 161 472 162 473
rect 162 472 163 473
rect 163 472 164 473
rect 214 472 215 473
rect 215 472 216 473
rect 216 472 217 473
rect 217 472 218 473
rect 218 472 219 473
rect 219 472 220 473
rect 220 472 221 473
rect 221 472 222 473
rect 222 472 223 473
rect 223 472 224 473
rect 224 472 225 473
rect 225 472 226 473
rect 226 472 227 473
rect 227 472 228 473
rect 228 472 229 473
rect 229 472 230 473
rect 230 472 231 473
rect 400 472 401 473
rect 401 472 402 473
rect 402 472 403 473
rect 403 472 404 473
rect 404 472 405 473
rect 405 472 406 473
rect 406 472 407 473
rect 407 472 408 473
rect 408 472 409 473
rect 409 472 410 473
rect 410 472 411 473
rect 411 472 412 473
rect 412 472 413 473
rect 413 472 414 473
rect 414 472 415 473
rect 137 471 138 472
rect 138 471 139 472
rect 139 471 140 472
rect 140 471 141 472
rect 141 471 142 472
rect 142 471 143 472
rect 143 471 144 472
rect 144 471 145 472
rect 145 471 146 472
rect 159 471 160 472
rect 160 471 161 472
rect 161 471 162 472
rect 162 471 163 472
rect 163 471 164 472
rect 164 471 165 472
rect 213 471 214 472
rect 214 471 215 472
rect 215 471 216 472
rect 216 471 217 472
rect 217 471 218 472
rect 218 471 219 472
rect 219 471 220 472
rect 220 471 221 472
rect 221 471 222 472
rect 222 471 223 472
rect 223 471 224 472
rect 224 471 225 472
rect 225 471 226 472
rect 226 471 227 472
rect 227 471 228 472
rect 228 471 229 472
rect 402 471 403 472
rect 403 471 404 472
rect 404 471 405 472
rect 405 471 406 472
rect 406 471 407 472
rect 407 471 408 472
rect 408 471 409 472
rect 409 471 410 472
rect 410 471 411 472
rect 411 471 412 472
rect 412 471 413 472
rect 413 471 414 472
rect 414 471 415 472
rect 415 471 416 472
rect 137 470 138 471
rect 138 470 139 471
rect 139 470 140 471
rect 140 470 141 471
rect 141 470 142 471
rect 142 470 143 471
rect 143 470 144 471
rect 144 470 145 471
rect 145 470 146 471
rect 146 470 147 471
rect 159 470 160 471
rect 160 470 161 471
rect 161 470 162 471
rect 162 470 163 471
rect 163 470 164 471
rect 164 470 165 471
rect 211 470 212 471
rect 212 470 213 471
rect 213 470 214 471
rect 214 470 215 471
rect 215 470 216 471
rect 216 470 217 471
rect 217 470 218 471
rect 218 470 219 471
rect 219 470 220 471
rect 220 470 221 471
rect 221 470 222 471
rect 222 470 223 471
rect 223 470 224 471
rect 224 470 225 471
rect 225 470 226 471
rect 226 470 227 471
rect 403 470 404 471
rect 404 470 405 471
rect 405 470 406 471
rect 406 470 407 471
rect 407 470 408 471
rect 408 470 409 471
rect 409 470 410 471
rect 410 470 411 471
rect 411 470 412 471
rect 412 470 413 471
rect 413 470 414 471
rect 414 470 415 471
rect 415 470 416 471
rect 416 470 417 471
rect 138 469 139 470
rect 139 469 140 470
rect 140 469 141 470
rect 141 469 142 470
rect 142 469 143 470
rect 143 469 144 470
rect 144 469 145 470
rect 145 469 146 470
rect 146 469 147 470
rect 159 469 160 470
rect 160 469 161 470
rect 161 469 162 470
rect 162 469 163 470
rect 163 469 164 470
rect 164 469 165 470
rect 210 469 211 470
rect 211 469 212 470
rect 212 469 213 470
rect 213 469 214 470
rect 214 469 215 470
rect 215 469 216 470
rect 216 469 217 470
rect 217 469 218 470
rect 218 469 219 470
rect 219 469 220 470
rect 220 469 221 470
rect 221 469 222 470
rect 222 469 223 470
rect 223 469 224 470
rect 224 469 225 470
rect 225 469 226 470
rect 404 469 405 470
rect 405 469 406 470
rect 406 469 407 470
rect 407 469 408 470
rect 408 469 409 470
rect 409 469 410 470
rect 410 469 411 470
rect 411 469 412 470
rect 412 469 413 470
rect 413 469 414 470
rect 414 469 415 470
rect 415 469 416 470
rect 416 469 417 470
rect 417 469 418 470
rect 418 469 419 470
rect 138 468 139 469
rect 139 468 140 469
rect 140 468 141 469
rect 141 468 142 469
rect 142 468 143 469
rect 143 468 144 469
rect 144 468 145 469
rect 145 468 146 469
rect 146 468 147 469
rect 160 468 161 469
rect 161 468 162 469
rect 162 468 163 469
rect 163 468 164 469
rect 164 468 165 469
rect 165 468 166 469
rect 208 468 209 469
rect 209 468 210 469
rect 210 468 211 469
rect 211 468 212 469
rect 212 468 213 469
rect 213 468 214 469
rect 214 468 215 469
rect 215 468 216 469
rect 216 468 217 469
rect 217 468 218 469
rect 218 468 219 469
rect 219 468 220 469
rect 220 468 221 469
rect 221 468 222 469
rect 222 468 223 469
rect 223 468 224 469
rect 406 468 407 469
rect 407 468 408 469
rect 408 468 409 469
rect 409 468 410 469
rect 410 468 411 469
rect 411 468 412 469
rect 412 468 413 469
rect 413 468 414 469
rect 414 468 415 469
rect 415 468 416 469
rect 416 468 417 469
rect 417 468 418 469
rect 418 468 419 469
rect 419 468 420 469
rect 138 467 139 468
rect 139 467 140 468
rect 140 467 141 468
rect 141 467 142 468
rect 142 467 143 468
rect 143 467 144 468
rect 144 467 145 468
rect 145 467 146 468
rect 146 467 147 468
rect 160 467 161 468
rect 161 467 162 468
rect 162 467 163 468
rect 163 467 164 468
rect 164 467 165 468
rect 165 467 166 468
rect 207 467 208 468
rect 208 467 209 468
rect 209 467 210 468
rect 210 467 211 468
rect 211 467 212 468
rect 212 467 213 468
rect 213 467 214 468
rect 214 467 215 468
rect 215 467 216 468
rect 216 467 217 468
rect 217 467 218 468
rect 218 467 219 468
rect 219 467 220 468
rect 220 467 221 468
rect 221 467 222 468
rect 407 467 408 468
rect 408 467 409 468
rect 409 467 410 468
rect 410 467 411 468
rect 411 467 412 468
rect 412 467 413 468
rect 413 467 414 468
rect 414 467 415 468
rect 415 467 416 468
rect 416 467 417 468
rect 417 467 418 468
rect 418 467 419 468
rect 419 467 420 468
rect 420 467 421 468
rect 139 466 140 467
rect 140 466 141 467
rect 141 466 142 467
rect 142 466 143 467
rect 143 466 144 467
rect 144 466 145 467
rect 145 466 146 467
rect 146 466 147 467
rect 147 466 148 467
rect 160 466 161 467
rect 161 466 162 467
rect 162 466 163 467
rect 163 466 164 467
rect 164 466 165 467
rect 165 466 166 467
rect 205 466 206 467
rect 206 466 207 467
rect 207 466 208 467
rect 208 466 209 467
rect 209 466 210 467
rect 210 466 211 467
rect 211 466 212 467
rect 212 466 213 467
rect 213 466 214 467
rect 214 466 215 467
rect 215 466 216 467
rect 216 466 217 467
rect 217 466 218 467
rect 218 466 219 467
rect 219 466 220 467
rect 220 466 221 467
rect 409 466 410 467
rect 410 466 411 467
rect 411 466 412 467
rect 412 466 413 467
rect 413 466 414 467
rect 414 466 415 467
rect 415 466 416 467
rect 416 466 417 467
rect 417 466 418 467
rect 418 466 419 467
rect 419 466 420 467
rect 420 466 421 467
rect 421 466 422 467
rect 422 466 423 467
rect 139 465 140 466
rect 140 465 141 466
rect 141 465 142 466
rect 142 465 143 466
rect 143 465 144 466
rect 144 465 145 466
rect 145 465 146 466
rect 146 465 147 466
rect 147 465 148 466
rect 160 465 161 466
rect 161 465 162 466
rect 162 465 163 466
rect 163 465 164 466
rect 164 465 165 466
rect 165 465 166 466
rect 204 465 205 466
rect 205 465 206 466
rect 206 465 207 466
rect 207 465 208 466
rect 208 465 209 466
rect 209 465 210 466
rect 210 465 211 466
rect 211 465 212 466
rect 212 465 213 466
rect 213 465 214 466
rect 214 465 215 466
rect 215 465 216 466
rect 216 465 217 466
rect 217 465 218 466
rect 218 465 219 466
rect 410 465 411 466
rect 411 465 412 466
rect 412 465 413 466
rect 413 465 414 466
rect 414 465 415 466
rect 415 465 416 466
rect 416 465 417 466
rect 417 465 418 466
rect 418 465 419 466
rect 419 465 420 466
rect 420 465 421 466
rect 421 465 422 466
rect 422 465 423 466
rect 423 465 424 466
rect 139 464 140 465
rect 140 464 141 465
rect 141 464 142 465
rect 142 464 143 465
rect 143 464 144 465
rect 144 464 145 465
rect 145 464 146 465
rect 146 464 147 465
rect 147 464 148 465
rect 161 464 162 465
rect 162 464 163 465
rect 163 464 164 465
rect 164 464 165 465
rect 165 464 166 465
rect 202 464 203 465
rect 203 464 204 465
rect 204 464 205 465
rect 205 464 206 465
rect 206 464 207 465
rect 207 464 208 465
rect 208 464 209 465
rect 209 464 210 465
rect 210 464 211 465
rect 211 464 212 465
rect 212 464 213 465
rect 213 464 214 465
rect 214 464 215 465
rect 215 464 216 465
rect 216 464 217 465
rect 411 464 412 465
rect 412 464 413 465
rect 413 464 414 465
rect 414 464 415 465
rect 415 464 416 465
rect 416 464 417 465
rect 417 464 418 465
rect 418 464 419 465
rect 419 464 420 465
rect 420 464 421 465
rect 421 464 422 465
rect 422 464 423 465
rect 423 464 424 465
rect 424 464 425 465
rect 139 463 140 464
rect 140 463 141 464
rect 141 463 142 464
rect 142 463 143 464
rect 143 463 144 464
rect 144 463 145 464
rect 145 463 146 464
rect 146 463 147 464
rect 147 463 148 464
rect 148 463 149 464
rect 161 463 162 464
rect 162 463 163 464
rect 163 463 164 464
rect 164 463 165 464
rect 165 463 166 464
rect 201 463 202 464
rect 202 463 203 464
rect 203 463 204 464
rect 204 463 205 464
rect 205 463 206 464
rect 206 463 207 464
rect 207 463 208 464
rect 208 463 209 464
rect 209 463 210 464
rect 210 463 211 464
rect 211 463 212 464
rect 212 463 213 464
rect 213 463 214 464
rect 214 463 215 464
rect 215 463 216 464
rect 413 463 414 464
rect 414 463 415 464
rect 415 463 416 464
rect 416 463 417 464
rect 417 463 418 464
rect 418 463 419 464
rect 419 463 420 464
rect 420 463 421 464
rect 421 463 422 464
rect 422 463 423 464
rect 423 463 424 464
rect 424 463 425 464
rect 425 463 426 464
rect 140 462 141 463
rect 141 462 142 463
rect 142 462 143 463
rect 143 462 144 463
rect 144 462 145 463
rect 145 462 146 463
rect 146 462 147 463
rect 147 462 148 463
rect 148 462 149 463
rect 161 462 162 463
rect 162 462 163 463
rect 163 462 164 463
rect 164 462 165 463
rect 165 462 166 463
rect 199 462 200 463
rect 200 462 201 463
rect 201 462 202 463
rect 202 462 203 463
rect 203 462 204 463
rect 204 462 205 463
rect 205 462 206 463
rect 206 462 207 463
rect 207 462 208 463
rect 208 462 209 463
rect 209 462 210 463
rect 210 462 211 463
rect 211 462 212 463
rect 212 462 213 463
rect 213 462 214 463
rect 414 462 415 463
rect 415 462 416 463
rect 416 462 417 463
rect 417 462 418 463
rect 418 462 419 463
rect 419 462 420 463
rect 420 462 421 463
rect 421 462 422 463
rect 422 462 423 463
rect 423 462 424 463
rect 424 462 425 463
rect 425 462 426 463
rect 426 462 427 463
rect 427 462 428 463
rect 140 461 141 462
rect 141 461 142 462
rect 142 461 143 462
rect 143 461 144 462
rect 144 461 145 462
rect 145 461 146 462
rect 146 461 147 462
rect 147 461 148 462
rect 148 461 149 462
rect 161 461 162 462
rect 162 461 163 462
rect 163 461 164 462
rect 164 461 165 462
rect 198 461 199 462
rect 199 461 200 462
rect 200 461 201 462
rect 201 461 202 462
rect 202 461 203 462
rect 203 461 204 462
rect 204 461 205 462
rect 205 461 206 462
rect 206 461 207 462
rect 207 461 208 462
rect 208 461 209 462
rect 209 461 210 462
rect 210 461 211 462
rect 211 461 212 462
rect 212 461 213 462
rect 415 461 416 462
rect 416 461 417 462
rect 417 461 418 462
rect 418 461 419 462
rect 419 461 420 462
rect 420 461 421 462
rect 421 461 422 462
rect 422 461 423 462
rect 423 461 424 462
rect 424 461 425 462
rect 425 461 426 462
rect 426 461 427 462
rect 427 461 428 462
rect 428 461 429 462
rect 140 460 141 461
rect 141 460 142 461
rect 142 460 143 461
rect 143 460 144 461
rect 144 460 145 461
rect 145 460 146 461
rect 146 460 147 461
rect 147 460 148 461
rect 148 460 149 461
rect 161 460 162 461
rect 162 460 163 461
rect 163 460 164 461
rect 197 460 198 461
rect 198 460 199 461
rect 199 460 200 461
rect 200 460 201 461
rect 201 460 202 461
rect 202 460 203 461
rect 203 460 204 461
rect 204 460 205 461
rect 205 460 206 461
rect 206 460 207 461
rect 207 460 208 461
rect 208 460 209 461
rect 209 460 210 461
rect 210 460 211 461
rect 417 460 418 461
rect 418 460 419 461
rect 419 460 420 461
rect 420 460 421 461
rect 421 460 422 461
rect 422 460 423 461
rect 423 460 424 461
rect 424 460 425 461
rect 425 460 426 461
rect 426 460 427 461
rect 427 460 428 461
rect 428 460 429 461
rect 429 460 430 461
rect 141 459 142 460
rect 142 459 143 460
rect 143 459 144 460
rect 144 459 145 460
rect 145 459 146 460
rect 146 459 147 460
rect 147 459 148 460
rect 148 459 149 460
rect 149 459 150 460
rect 195 459 196 460
rect 196 459 197 460
rect 197 459 198 460
rect 198 459 199 460
rect 199 459 200 460
rect 200 459 201 460
rect 201 459 202 460
rect 202 459 203 460
rect 203 459 204 460
rect 204 459 205 460
rect 205 459 206 460
rect 206 459 207 460
rect 207 459 208 460
rect 208 459 209 460
rect 209 459 210 460
rect 418 459 419 460
rect 419 459 420 460
rect 420 459 421 460
rect 421 459 422 460
rect 422 459 423 460
rect 423 459 424 460
rect 424 459 425 460
rect 425 459 426 460
rect 426 459 427 460
rect 427 459 428 460
rect 428 459 429 460
rect 429 459 430 460
rect 430 459 431 460
rect 431 459 432 460
rect 141 458 142 459
rect 142 458 143 459
rect 143 458 144 459
rect 144 458 145 459
rect 145 458 146 459
rect 146 458 147 459
rect 147 458 148 459
rect 148 458 149 459
rect 149 458 150 459
rect 194 458 195 459
rect 195 458 196 459
rect 196 458 197 459
rect 197 458 198 459
rect 198 458 199 459
rect 199 458 200 459
rect 200 458 201 459
rect 201 458 202 459
rect 202 458 203 459
rect 203 458 204 459
rect 204 458 205 459
rect 205 458 206 459
rect 206 458 207 459
rect 207 458 208 459
rect 419 458 420 459
rect 420 458 421 459
rect 421 458 422 459
rect 422 458 423 459
rect 423 458 424 459
rect 424 458 425 459
rect 425 458 426 459
rect 426 458 427 459
rect 427 458 428 459
rect 428 458 429 459
rect 429 458 430 459
rect 430 458 431 459
rect 431 458 432 459
rect 432 458 433 459
rect 141 457 142 458
rect 142 457 143 458
rect 143 457 144 458
rect 144 457 145 458
rect 145 457 146 458
rect 146 457 147 458
rect 147 457 148 458
rect 148 457 149 458
rect 149 457 150 458
rect 193 457 194 458
rect 194 457 195 458
rect 195 457 196 458
rect 196 457 197 458
rect 197 457 198 458
rect 198 457 199 458
rect 199 457 200 458
rect 200 457 201 458
rect 201 457 202 458
rect 202 457 203 458
rect 203 457 204 458
rect 204 457 205 458
rect 205 457 206 458
rect 206 457 207 458
rect 421 457 422 458
rect 422 457 423 458
rect 423 457 424 458
rect 424 457 425 458
rect 425 457 426 458
rect 426 457 427 458
rect 427 457 428 458
rect 428 457 429 458
rect 429 457 430 458
rect 430 457 431 458
rect 431 457 432 458
rect 432 457 433 458
rect 433 457 434 458
rect 141 456 142 457
rect 142 456 143 457
rect 143 456 144 457
rect 144 456 145 457
rect 145 456 146 457
rect 146 456 147 457
rect 147 456 148 457
rect 148 456 149 457
rect 149 456 150 457
rect 150 456 151 457
rect 191 456 192 457
rect 192 456 193 457
rect 193 456 194 457
rect 194 456 195 457
rect 195 456 196 457
rect 196 456 197 457
rect 197 456 198 457
rect 198 456 199 457
rect 199 456 200 457
rect 200 456 201 457
rect 201 456 202 457
rect 202 456 203 457
rect 203 456 204 457
rect 204 456 205 457
rect 422 456 423 457
rect 423 456 424 457
rect 424 456 425 457
rect 425 456 426 457
rect 426 456 427 457
rect 427 456 428 457
rect 428 456 429 457
rect 429 456 430 457
rect 430 456 431 457
rect 431 456 432 457
rect 432 456 433 457
rect 433 456 434 457
rect 434 456 435 457
rect 142 455 143 456
rect 143 455 144 456
rect 144 455 145 456
rect 145 455 146 456
rect 146 455 147 456
rect 147 455 148 456
rect 148 455 149 456
rect 149 455 150 456
rect 150 455 151 456
rect 190 455 191 456
rect 191 455 192 456
rect 192 455 193 456
rect 193 455 194 456
rect 194 455 195 456
rect 195 455 196 456
rect 196 455 197 456
rect 197 455 198 456
rect 198 455 199 456
rect 199 455 200 456
rect 200 455 201 456
rect 201 455 202 456
rect 202 455 203 456
rect 203 455 204 456
rect 423 455 424 456
rect 424 455 425 456
rect 425 455 426 456
rect 426 455 427 456
rect 427 455 428 456
rect 428 455 429 456
rect 429 455 430 456
rect 430 455 431 456
rect 431 455 432 456
rect 432 455 433 456
rect 433 455 434 456
rect 434 455 435 456
rect 435 455 436 456
rect 142 454 143 455
rect 143 454 144 455
rect 144 454 145 455
rect 145 454 146 455
rect 146 454 147 455
rect 147 454 148 455
rect 148 454 149 455
rect 149 454 150 455
rect 150 454 151 455
rect 189 454 190 455
rect 190 454 191 455
rect 191 454 192 455
rect 192 454 193 455
rect 193 454 194 455
rect 194 454 195 455
rect 195 454 196 455
rect 196 454 197 455
rect 197 454 198 455
rect 198 454 199 455
rect 199 454 200 455
rect 200 454 201 455
rect 201 454 202 455
rect 202 454 203 455
rect 425 454 426 455
rect 426 454 427 455
rect 427 454 428 455
rect 428 454 429 455
rect 429 454 430 455
rect 430 454 431 455
rect 431 454 432 455
rect 432 454 433 455
rect 433 454 434 455
rect 434 454 435 455
rect 435 454 436 455
rect 436 454 437 455
rect 437 454 438 455
rect 142 453 143 454
rect 143 453 144 454
rect 144 453 145 454
rect 145 453 146 454
rect 146 453 147 454
rect 147 453 148 454
rect 148 453 149 454
rect 149 453 150 454
rect 150 453 151 454
rect 187 453 188 454
rect 188 453 189 454
rect 189 453 190 454
rect 190 453 191 454
rect 191 453 192 454
rect 192 453 193 454
rect 193 453 194 454
rect 194 453 195 454
rect 195 453 196 454
rect 196 453 197 454
rect 197 453 198 454
rect 198 453 199 454
rect 199 453 200 454
rect 200 453 201 454
rect 426 453 427 454
rect 427 453 428 454
rect 428 453 429 454
rect 429 453 430 454
rect 430 453 431 454
rect 431 453 432 454
rect 432 453 433 454
rect 433 453 434 454
rect 434 453 435 454
rect 435 453 436 454
rect 436 453 437 454
rect 437 453 438 454
rect 438 453 439 454
rect 142 452 143 453
rect 143 452 144 453
rect 144 452 145 453
rect 145 452 146 453
rect 146 452 147 453
rect 147 452 148 453
rect 148 452 149 453
rect 149 452 150 453
rect 150 452 151 453
rect 151 452 152 453
rect 186 452 187 453
rect 187 452 188 453
rect 188 452 189 453
rect 189 452 190 453
rect 190 452 191 453
rect 191 452 192 453
rect 192 452 193 453
rect 193 452 194 453
rect 194 452 195 453
rect 195 452 196 453
rect 196 452 197 453
rect 197 452 198 453
rect 198 452 199 453
rect 199 452 200 453
rect 427 452 428 453
rect 428 452 429 453
rect 429 452 430 453
rect 430 452 431 453
rect 431 452 432 453
rect 432 452 433 453
rect 433 452 434 453
rect 434 452 435 453
rect 435 452 436 453
rect 436 452 437 453
rect 437 452 438 453
rect 438 452 439 453
rect 439 452 440 453
rect 143 451 144 452
rect 144 451 145 452
rect 145 451 146 452
rect 146 451 147 452
rect 147 451 148 452
rect 148 451 149 452
rect 149 451 150 452
rect 150 451 151 452
rect 151 451 152 452
rect 185 451 186 452
rect 186 451 187 452
rect 187 451 188 452
rect 188 451 189 452
rect 189 451 190 452
rect 190 451 191 452
rect 191 451 192 452
rect 192 451 193 452
rect 193 451 194 452
rect 194 451 195 452
rect 195 451 196 452
rect 196 451 197 452
rect 197 451 198 452
rect 198 451 199 452
rect 428 451 429 452
rect 429 451 430 452
rect 430 451 431 452
rect 431 451 432 452
rect 432 451 433 452
rect 433 451 434 452
rect 434 451 435 452
rect 435 451 436 452
rect 436 451 437 452
rect 437 451 438 452
rect 438 451 439 452
rect 439 451 440 452
rect 440 451 441 452
rect 143 450 144 451
rect 144 450 145 451
rect 145 450 146 451
rect 146 450 147 451
rect 147 450 148 451
rect 148 450 149 451
rect 149 450 150 451
rect 150 450 151 451
rect 151 450 152 451
rect 184 450 185 451
rect 185 450 186 451
rect 186 450 187 451
rect 187 450 188 451
rect 188 450 189 451
rect 189 450 190 451
rect 190 450 191 451
rect 191 450 192 451
rect 192 450 193 451
rect 193 450 194 451
rect 194 450 195 451
rect 195 450 196 451
rect 196 450 197 451
rect 429 450 430 451
rect 430 450 431 451
rect 431 450 432 451
rect 432 450 433 451
rect 433 450 434 451
rect 434 450 435 451
rect 435 450 436 451
rect 436 450 437 451
rect 437 450 438 451
rect 438 450 439 451
rect 439 450 440 451
rect 440 450 441 451
rect 441 450 442 451
rect 143 449 144 450
rect 144 449 145 450
rect 145 449 146 450
rect 146 449 147 450
rect 147 449 148 450
rect 148 449 149 450
rect 149 449 150 450
rect 150 449 151 450
rect 151 449 152 450
rect 183 449 184 450
rect 184 449 185 450
rect 185 449 186 450
rect 186 449 187 450
rect 187 449 188 450
rect 188 449 189 450
rect 189 449 190 450
rect 190 449 191 450
rect 191 449 192 450
rect 192 449 193 450
rect 193 449 194 450
rect 194 449 195 450
rect 195 449 196 450
rect 431 449 432 450
rect 432 449 433 450
rect 433 449 434 450
rect 434 449 435 450
rect 435 449 436 450
rect 436 449 437 450
rect 437 449 438 450
rect 438 449 439 450
rect 439 449 440 450
rect 440 449 441 450
rect 441 449 442 450
rect 442 449 443 450
rect 143 448 144 449
rect 144 448 145 449
rect 145 448 146 449
rect 146 448 147 449
rect 147 448 148 449
rect 148 448 149 449
rect 149 448 150 449
rect 150 448 151 449
rect 151 448 152 449
rect 152 448 153 449
rect 181 448 182 449
rect 182 448 183 449
rect 183 448 184 449
rect 184 448 185 449
rect 185 448 186 449
rect 186 448 187 449
rect 187 448 188 449
rect 188 448 189 449
rect 189 448 190 449
rect 190 448 191 449
rect 191 448 192 449
rect 192 448 193 449
rect 193 448 194 449
rect 194 448 195 449
rect 432 448 433 449
rect 433 448 434 449
rect 434 448 435 449
rect 435 448 436 449
rect 436 448 437 449
rect 437 448 438 449
rect 438 448 439 449
rect 439 448 440 449
rect 440 448 441 449
rect 441 448 442 449
rect 442 448 443 449
rect 443 448 444 449
rect 444 448 445 449
rect 144 447 145 448
rect 145 447 146 448
rect 146 447 147 448
rect 147 447 148 448
rect 148 447 149 448
rect 149 447 150 448
rect 150 447 151 448
rect 151 447 152 448
rect 152 447 153 448
rect 180 447 181 448
rect 181 447 182 448
rect 182 447 183 448
rect 183 447 184 448
rect 184 447 185 448
rect 185 447 186 448
rect 186 447 187 448
rect 187 447 188 448
rect 188 447 189 448
rect 189 447 190 448
rect 190 447 191 448
rect 191 447 192 448
rect 192 447 193 448
rect 433 447 434 448
rect 434 447 435 448
rect 435 447 436 448
rect 436 447 437 448
rect 437 447 438 448
rect 438 447 439 448
rect 439 447 440 448
rect 440 447 441 448
rect 441 447 442 448
rect 442 447 443 448
rect 443 447 444 448
rect 444 447 445 448
rect 445 447 446 448
rect 144 446 145 447
rect 145 446 146 447
rect 146 446 147 447
rect 147 446 148 447
rect 148 446 149 447
rect 149 446 150 447
rect 150 446 151 447
rect 151 446 152 447
rect 152 446 153 447
rect 179 446 180 447
rect 180 446 181 447
rect 181 446 182 447
rect 182 446 183 447
rect 183 446 184 447
rect 184 446 185 447
rect 185 446 186 447
rect 186 446 187 447
rect 187 446 188 447
rect 188 446 189 447
rect 189 446 190 447
rect 190 446 191 447
rect 191 446 192 447
rect 434 446 435 447
rect 435 446 436 447
rect 436 446 437 447
rect 437 446 438 447
rect 438 446 439 447
rect 439 446 440 447
rect 440 446 441 447
rect 441 446 442 447
rect 442 446 443 447
rect 443 446 444 447
rect 444 446 445 447
rect 445 446 446 447
rect 446 446 447 447
rect 144 445 145 446
rect 145 445 146 446
rect 146 445 147 446
rect 147 445 148 446
rect 148 445 149 446
rect 149 445 150 446
rect 150 445 151 446
rect 151 445 152 446
rect 152 445 153 446
rect 178 445 179 446
rect 179 445 180 446
rect 180 445 181 446
rect 181 445 182 446
rect 182 445 183 446
rect 183 445 184 446
rect 184 445 185 446
rect 185 445 186 446
rect 186 445 187 446
rect 187 445 188 446
rect 188 445 189 446
rect 189 445 190 446
rect 190 445 191 446
rect 435 445 436 446
rect 436 445 437 446
rect 437 445 438 446
rect 438 445 439 446
rect 439 445 440 446
rect 440 445 441 446
rect 441 445 442 446
rect 442 445 443 446
rect 443 445 444 446
rect 444 445 445 446
rect 445 445 446 446
rect 446 445 447 446
rect 447 445 448 446
rect 144 444 145 445
rect 145 444 146 445
rect 146 444 147 445
rect 147 444 148 445
rect 148 444 149 445
rect 149 444 150 445
rect 150 444 151 445
rect 151 444 152 445
rect 152 444 153 445
rect 153 444 154 445
rect 177 444 178 445
rect 178 444 179 445
rect 179 444 180 445
rect 180 444 181 445
rect 181 444 182 445
rect 182 444 183 445
rect 183 444 184 445
rect 184 444 185 445
rect 185 444 186 445
rect 186 444 187 445
rect 187 444 188 445
rect 188 444 189 445
rect 189 444 190 445
rect 437 444 438 445
rect 438 444 439 445
rect 439 444 440 445
rect 440 444 441 445
rect 441 444 442 445
rect 442 444 443 445
rect 443 444 444 445
rect 444 444 445 445
rect 445 444 446 445
rect 446 444 447 445
rect 447 444 448 445
rect 448 444 449 445
rect 145 443 146 444
rect 146 443 147 444
rect 147 443 148 444
rect 148 443 149 444
rect 149 443 150 444
rect 150 443 151 444
rect 151 443 152 444
rect 152 443 153 444
rect 153 443 154 444
rect 176 443 177 444
rect 177 443 178 444
rect 178 443 179 444
rect 179 443 180 444
rect 180 443 181 444
rect 181 443 182 444
rect 182 443 183 444
rect 183 443 184 444
rect 184 443 185 444
rect 185 443 186 444
rect 186 443 187 444
rect 187 443 188 444
rect 188 443 189 444
rect 438 443 439 444
rect 439 443 440 444
rect 440 443 441 444
rect 441 443 442 444
rect 442 443 443 444
rect 443 443 444 444
rect 444 443 445 444
rect 445 443 446 444
rect 446 443 447 444
rect 447 443 448 444
rect 448 443 449 444
rect 449 443 450 444
rect 145 442 146 443
rect 146 442 147 443
rect 147 442 148 443
rect 148 442 149 443
rect 149 442 150 443
rect 150 442 151 443
rect 151 442 152 443
rect 152 442 153 443
rect 153 442 154 443
rect 175 442 176 443
rect 176 442 177 443
rect 177 442 178 443
rect 178 442 179 443
rect 179 442 180 443
rect 180 442 181 443
rect 181 442 182 443
rect 182 442 183 443
rect 183 442 184 443
rect 184 442 185 443
rect 185 442 186 443
rect 186 442 187 443
rect 439 442 440 443
rect 440 442 441 443
rect 441 442 442 443
rect 442 442 443 443
rect 443 442 444 443
rect 444 442 445 443
rect 445 442 446 443
rect 446 442 447 443
rect 447 442 448 443
rect 448 442 449 443
rect 449 442 450 443
rect 450 442 451 443
rect 145 441 146 442
rect 146 441 147 442
rect 147 441 148 442
rect 148 441 149 442
rect 149 441 150 442
rect 150 441 151 442
rect 151 441 152 442
rect 152 441 153 442
rect 153 441 154 442
rect 174 441 175 442
rect 175 441 176 442
rect 176 441 177 442
rect 177 441 178 442
rect 178 441 179 442
rect 179 441 180 442
rect 180 441 181 442
rect 181 441 182 442
rect 182 441 183 442
rect 183 441 184 442
rect 184 441 185 442
rect 185 441 186 442
rect 440 441 441 442
rect 441 441 442 442
rect 442 441 443 442
rect 443 441 444 442
rect 444 441 445 442
rect 445 441 446 442
rect 446 441 447 442
rect 447 441 448 442
rect 448 441 449 442
rect 449 441 450 442
rect 450 441 451 442
rect 451 441 452 442
rect 145 440 146 441
rect 146 440 147 441
rect 147 440 148 441
rect 148 440 149 441
rect 149 440 150 441
rect 150 440 151 441
rect 151 440 152 441
rect 152 440 153 441
rect 153 440 154 441
rect 173 440 174 441
rect 174 440 175 441
rect 175 440 176 441
rect 176 440 177 441
rect 177 440 178 441
rect 178 440 179 441
rect 179 440 180 441
rect 180 440 181 441
rect 181 440 182 441
rect 182 440 183 441
rect 183 440 184 441
rect 184 440 185 441
rect 441 440 442 441
rect 442 440 443 441
rect 443 440 444 441
rect 444 440 445 441
rect 445 440 446 441
rect 446 440 447 441
rect 447 440 448 441
rect 448 440 449 441
rect 449 440 450 441
rect 450 440 451 441
rect 451 440 452 441
rect 452 440 453 441
rect 146 439 147 440
rect 147 439 148 440
rect 148 439 149 440
rect 149 439 150 440
rect 150 439 151 440
rect 151 439 152 440
rect 152 439 153 440
rect 153 439 154 440
rect 154 439 155 440
rect 172 439 173 440
rect 173 439 174 440
rect 174 439 175 440
rect 175 439 176 440
rect 176 439 177 440
rect 177 439 178 440
rect 178 439 179 440
rect 179 439 180 440
rect 180 439 181 440
rect 181 439 182 440
rect 182 439 183 440
rect 183 439 184 440
rect 442 439 443 440
rect 443 439 444 440
rect 444 439 445 440
rect 445 439 446 440
rect 446 439 447 440
rect 447 439 448 440
rect 448 439 449 440
rect 449 439 450 440
rect 450 439 451 440
rect 451 439 452 440
rect 452 439 453 440
rect 453 439 454 440
rect 454 439 455 440
rect 146 438 147 439
rect 147 438 148 439
rect 148 438 149 439
rect 149 438 150 439
rect 150 438 151 439
rect 151 438 152 439
rect 152 438 153 439
rect 153 438 154 439
rect 154 438 155 439
rect 171 438 172 439
rect 172 438 173 439
rect 173 438 174 439
rect 174 438 175 439
rect 175 438 176 439
rect 176 438 177 439
rect 177 438 178 439
rect 178 438 179 439
rect 179 438 180 439
rect 180 438 181 439
rect 181 438 182 439
rect 182 438 183 439
rect 443 438 444 439
rect 444 438 445 439
rect 445 438 446 439
rect 446 438 447 439
rect 447 438 448 439
rect 448 438 449 439
rect 449 438 450 439
rect 450 438 451 439
rect 451 438 452 439
rect 452 438 453 439
rect 453 438 454 439
rect 454 438 455 439
rect 455 438 456 439
rect 146 437 147 438
rect 147 437 148 438
rect 148 437 149 438
rect 149 437 150 438
rect 150 437 151 438
rect 151 437 152 438
rect 152 437 153 438
rect 153 437 154 438
rect 154 437 155 438
rect 170 437 171 438
rect 171 437 172 438
rect 172 437 173 438
rect 173 437 174 438
rect 174 437 175 438
rect 175 437 176 438
rect 176 437 177 438
rect 177 437 178 438
rect 178 437 179 438
rect 179 437 180 438
rect 180 437 181 438
rect 181 437 182 438
rect 444 437 445 438
rect 445 437 446 438
rect 446 437 447 438
rect 447 437 448 438
rect 448 437 449 438
rect 449 437 450 438
rect 450 437 451 438
rect 451 437 452 438
rect 452 437 453 438
rect 453 437 454 438
rect 454 437 455 438
rect 455 437 456 438
rect 456 437 457 438
rect 146 436 147 437
rect 147 436 148 437
rect 148 436 149 437
rect 149 436 150 437
rect 150 436 151 437
rect 151 436 152 437
rect 152 436 153 437
rect 153 436 154 437
rect 154 436 155 437
rect 169 436 170 437
rect 170 436 171 437
rect 171 436 172 437
rect 172 436 173 437
rect 173 436 174 437
rect 174 436 175 437
rect 175 436 176 437
rect 176 436 177 437
rect 177 436 178 437
rect 178 436 179 437
rect 179 436 180 437
rect 180 436 181 437
rect 446 436 447 437
rect 447 436 448 437
rect 448 436 449 437
rect 449 436 450 437
rect 450 436 451 437
rect 451 436 452 437
rect 452 436 453 437
rect 453 436 454 437
rect 454 436 455 437
rect 455 436 456 437
rect 456 436 457 437
rect 457 436 458 437
rect 147 435 148 436
rect 148 435 149 436
rect 149 435 150 436
rect 150 435 151 436
rect 151 435 152 436
rect 152 435 153 436
rect 153 435 154 436
rect 154 435 155 436
rect 155 435 156 436
rect 168 435 169 436
rect 169 435 170 436
rect 170 435 171 436
rect 171 435 172 436
rect 172 435 173 436
rect 173 435 174 436
rect 174 435 175 436
rect 175 435 176 436
rect 176 435 177 436
rect 177 435 178 436
rect 178 435 179 436
rect 179 435 180 436
rect 447 435 448 436
rect 448 435 449 436
rect 449 435 450 436
rect 450 435 451 436
rect 451 435 452 436
rect 452 435 453 436
rect 453 435 454 436
rect 454 435 455 436
rect 455 435 456 436
rect 456 435 457 436
rect 457 435 458 436
rect 458 435 459 436
rect 147 434 148 435
rect 148 434 149 435
rect 149 434 150 435
rect 150 434 151 435
rect 151 434 152 435
rect 152 434 153 435
rect 153 434 154 435
rect 154 434 155 435
rect 155 434 156 435
rect 167 434 168 435
rect 168 434 169 435
rect 169 434 170 435
rect 170 434 171 435
rect 171 434 172 435
rect 172 434 173 435
rect 173 434 174 435
rect 174 434 175 435
rect 175 434 176 435
rect 176 434 177 435
rect 177 434 178 435
rect 178 434 179 435
rect 448 434 449 435
rect 449 434 450 435
rect 450 434 451 435
rect 451 434 452 435
rect 452 434 453 435
rect 453 434 454 435
rect 454 434 455 435
rect 455 434 456 435
rect 456 434 457 435
rect 457 434 458 435
rect 458 434 459 435
rect 459 434 460 435
rect 147 433 148 434
rect 148 433 149 434
rect 149 433 150 434
rect 150 433 151 434
rect 151 433 152 434
rect 152 433 153 434
rect 153 433 154 434
rect 154 433 155 434
rect 155 433 156 434
rect 166 433 167 434
rect 167 433 168 434
rect 168 433 169 434
rect 169 433 170 434
rect 170 433 171 434
rect 171 433 172 434
rect 172 433 173 434
rect 173 433 174 434
rect 174 433 175 434
rect 175 433 176 434
rect 176 433 177 434
rect 177 433 178 434
rect 449 433 450 434
rect 450 433 451 434
rect 451 433 452 434
rect 452 433 453 434
rect 453 433 454 434
rect 454 433 455 434
rect 455 433 456 434
rect 456 433 457 434
rect 457 433 458 434
rect 458 433 459 434
rect 459 433 460 434
rect 460 433 461 434
rect 147 432 148 433
rect 148 432 149 433
rect 149 432 150 433
rect 150 432 151 433
rect 151 432 152 433
rect 152 432 153 433
rect 153 432 154 433
rect 154 432 155 433
rect 155 432 156 433
rect 165 432 166 433
rect 166 432 167 433
rect 167 432 168 433
rect 168 432 169 433
rect 169 432 170 433
rect 170 432 171 433
rect 171 432 172 433
rect 172 432 173 433
rect 173 432 174 433
rect 174 432 175 433
rect 175 432 176 433
rect 176 432 177 433
rect 450 432 451 433
rect 451 432 452 433
rect 452 432 453 433
rect 453 432 454 433
rect 454 432 455 433
rect 455 432 456 433
rect 456 432 457 433
rect 457 432 458 433
rect 458 432 459 433
rect 459 432 460 433
rect 460 432 461 433
rect 461 432 462 433
rect 148 431 149 432
rect 149 431 150 432
rect 150 431 151 432
rect 151 431 152 432
rect 152 431 153 432
rect 153 431 154 432
rect 154 431 155 432
rect 155 431 156 432
rect 156 431 157 432
rect 164 431 165 432
rect 165 431 166 432
rect 166 431 167 432
rect 167 431 168 432
rect 168 431 169 432
rect 169 431 170 432
rect 170 431 171 432
rect 171 431 172 432
rect 172 431 173 432
rect 173 431 174 432
rect 174 431 175 432
rect 175 431 176 432
rect 451 431 452 432
rect 452 431 453 432
rect 453 431 454 432
rect 454 431 455 432
rect 455 431 456 432
rect 456 431 457 432
rect 457 431 458 432
rect 458 431 459 432
rect 459 431 460 432
rect 460 431 461 432
rect 461 431 462 432
rect 462 431 463 432
rect 148 430 149 431
rect 149 430 150 431
rect 150 430 151 431
rect 151 430 152 431
rect 152 430 153 431
rect 153 430 154 431
rect 154 430 155 431
rect 155 430 156 431
rect 156 430 157 431
rect 163 430 164 431
rect 164 430 165 431
rect 165 430 166 431
rect 166 430 167 431
rect 167 430 168 431
rect 168 430 169 431
rect 169 430 170 431
rect 170 430 171 431
rect 171 430 172 431
rect 172 430 173 431
rect 173 430 174 431
rect 174 430 175 431
rect 452 430 453 431
rect 453 430 454 431
rect 454 430 455 431
rect 455 430 456 431
rect 456 430 457 431
rect 457 430 458 431
rect 458 430 459 431
rect 459 430 460 431
rect 460 430 461 431
rect 461 430 462 431
rect 462 430 463 431
rect 463 430 464 431
rect 148 429 149 430
rect 149 429 150 430
rect 150 429 151 430
rect 151 429 152 430
rect 152 429 153 430
rect 153 429 154 430
rect 154 429 155 430
rect 155 429 156 430
rect 156 429 157 430
rect 162 429 163 430
rect 163 429 164 430
rect 164 429 165 430
rect 165 429 166 430
rect 166 429 167 430
rect 167 429 168 430
rect 168 429 169 430
rect 169 429 170 430
rect 170 429 171 430
rect 171 429 172 430
rect 172 429 173 430
rect 173 429 174 430
rect 453 429 454 430
rect 454 429 455 430
rect 455 429 456 430
rect 456 429 457 430
rect 457 429 458 430
rect 458 429 459 430
rect 459 429 460 430
rect 460 429 461 430
rect 461 429 462 430
rect 462 429 463 430
rect 463 429 464 430
rect 464 429 465 430
rect 148 428 149 429
rect 149 428 150 429
rect 150 428 151 429
rect 151 428 152 429
rect 152 428 153 429
rect 153 428 154 429
rect 154 428 155 429
rect 155 428 156 429
rect 156 428 157 429
rect 161 428 162 429
rect 162 428 163 429
rect 163 428 164 429
rect 164 428 165 429
rect 165 428 166 429
rect 166 428 167 429
rect 167 428 168 429
rect 168 428 169 429
rect 169 428 170 429
rect 170 428 171 429
rect 171 428 172 429
rect 172 428 173 429
rect 454 428 455 429
rect 455 428 456 429
rect 456 428 457 429
rect 457 428 458 429
rect 458 428 459 429
rect 459 428 460 429
rect 460 428 461 429
rect 461 428 462 429
rect 462 428 463 429
rect 463 428 464 429
rect 464 428 465 429
rect 465 428 466 429
rect 148 427 149 428
rect 149 427 150 428
rect 150 427 151 428
rect 151 427 152 428
rect 152 427 153 428
rect 153 427 154 428
rect 154 427 155 428
rect 155 427 156 428
rect 156 427 157 428
rect 160 427 161 428
rect 161 427 162 428
rect 162 427 163 428
rect 163 427 164 428
rect 164 427 165 428
rect 165 427 166 428
rect 166 427 167 428
rect 167 427 168 428
rect 168 427 169 428
rect 169 427 170 428
rect 170 427 171 428
rect 171 427 172 428
rect 455 427 456 428
rect 456 427 457 428
rect 457 427 458 428
rect 458 427 459 428
rect 459 427 460 428
rect 460 427 461 428
rect 461 427 462 428
rect 462 427 463 428
rect 463 427 464 428
rect 464 427 465 428
rect 465 427 466 428
rect 466 427 467 428
rect 149 426 150 427
rect 150 426 151 427
rect 151 426 152 427
rect 152 426 153 427
rect 153 426 154 427
rect 154 426 155 427
rect 155 426 156 427
rect 156 426 157 427
rect 157 426 158 427
rect 159 426 160 427
rect 160 426 161 427
rect 161 426 162 427
rect 162 426 163 427
rect 163 426 164 427
rect 164 426 165 427
rect 165 426 166 427
rect 166 426 167 427
rect 167 426 168 427
rect 168 426 169 427
rect 169 426 170 427
rect 170 426 171 427
rect 456 426 457 427
rect 457 426 458 427
rect 458 426 459 427
rect 459 426 460 427
rect 460 426 461 427
rect 461 426 462 427
rect 462 426 463 427
rect 463 426 464 427
rect 464 426 465 427
rect 465 426 466 427
rect 466 426 467 427
rect 467 426 468 427
rect 149 425 150 426
rect 150 425 151 426
rect 151 425 152 426
rect 152 425 153 426
rect 153 425 154 426
rect 154 425 155 426
rect 155 425 156 426
rect 156 425 157 426
rect 157 425 158 426
rect 158 425 159 426
rect 159 425 160 426
rect 160 425 161 426
rect 161 425 162 426
rect 162 425 163 426
rect 163 425 164 426
rect 164 425 165 426
rect 165 425 166 426
rect 166 425 167 426
rect 167 425 168 426
rect 168 425 169 426
rect 169 425 170 426
rect 457 425 458 426
rect 458 425 459 426
rect 459 425 460 426
rect 460 425 461 426
rect 461 425 462 426
rect 462 425 463 426
rect 463 425 464 426
rect 464 425 465 426
rect 465 425 466 426
rect 466 425 467 426
rect 467 425 468 426
rect 468 425 469 426
rect 149 424 150 425
rect 150 424 151 425
rect 151 424 152 425
rect 152 424 153 425
rect 153 424 154 425
rect 154 424 155 425
rect 155 424 156 425
rect 156 424 157 425
rect 157 424 158 425
rect 158 424 159 425
rect 159 424 160 425
rect 160 424 161 425
rect 161 424 162 425
rect 162 424 163 425
rect 163 424 164 425
rect 164 424 165 425
rect 165 424 166 425
rect 166 424 167 425
rect 167 424 168 425
rect 168 424 169 425
rect 458 424 459 425
rect 459 424 460 425
rect 460 424 461 425
rect 461 424 462 425
rect 462 424 463 425
rect 463 424 464 425
rect 464 424 465 425
rect 465 424 466 425
rect 466 424 467 425
rect 467 424 468 425
rect 468 424 469 425
rect 119 423 120 424
rect 120 423 121 424
rect 149 423 150 424
rect 150 423 151 424
rect 151 423 152 424
rect 152 423 153 424
rect 153 423 154 424
rect 154 423 155 424
rect 155 423 156 424
rect 156 423 157 424
rect 157 423 158 424
rect 158 423 159 424
rect 159 423 160 424
rect 160 423 161 424
rect 161 423 162 424
rect 162 423 163 424
rect 163 423 164 424
rect 164 423 165 424
rect 165 423 166 424
rect 166 423 167 424
rect 167 423 168 424
rect 459 423 460 424
rect 460 423 461 424
rect 461 423 462 424
rect 462 423 463 424
rect 463 423 464 424
rect 464 423 465 424
rect 465 423 466 424
rect 466 423 467 424
rect 467 423 468 424
rect 468 423 469 424
rect 469 423 470 424
rect 111 422 112 423
rect 112 422 113 423
rect 113 422 114 423
rect 114 422 115 423
rect 115 422 116 423
rect 116 422 117 423
rect 117 422 118 423
rect 118 422 119 423
rect 119 422 120 423
rect 120 422 121 423
rect 121 422 122 423
rect 122 422 123 423
rect 123 422 124 423
rect 124 422 125 423
rect 125 422 126 423
rect 126 422 127 423
rect 127 422 128 423
rect 128 422 129 423
rect 129 422 130 423
rect 130 422 131 423
rect 150 422 151 423
rect 151 422 152 423
rect 152 422 153 423
rect 153 422 154 423
rect 154 422 155 423
rect 155 422 156 423
rect 156 422 157 423
rect 157 422 158 423
rect 158 422 159 423
rect 159 422 160 423
rect 160 422 161 423
rect 161 422 162 423
rect 162 422 163 423
rect 163 422 164 423
rect 164 422 165 423
rect 165 422 166 423
rect 166 422 167 423
rect 460 422 461 423
rect 461 422 462 423
rect 462 422 463 423
rect 463 422 464 423
rect 464 422 465 423
rect 465 422 466 423
rect 466 422 467 423
rect 467 422 468 423
rect 468 422 469 423
rect 469 422 470 423
rect 470 422 471 423
rect 107 421 108 422
rect 108 421 109 422
rect 109 421 110 422
rect 110 421 111 422
rect 111 421 112 422
rect 112 421 113 422
rect 113 421 114 422
rect 114 421 115 422
rect 115 421 116 422
rect 116 421 117 422
rect 117 421 118 422
rect 118 421 119 422
rect 119 421 120 422
rect 120 421 121 422
rect 121 421 122 422
rect 122 421 123 422
rect 123 421 124 422
rect 124 421 125 422
rect 125 421 126 422
rect 126 421 127 422
rect 127 421 128 422
rect 128 421 129 422
rect 129 421 130 422
rect 130 421 131 422
rect 131 421 132 422
rect 132 421 133 422
rect 133 421 134 422
rect 134 421 135 422
rect 150 421 151 422
rect 151 421 152 422
rect 152 421 153 422
rect 153 421 154 422
rect 154 421 155 422
rect 155 421 156 422
rect 156 421 157 422
rect 157 421 158 422
rect 158 421 159 422
rect 159 421 160 422
rect 160 421 161 422
rect 161 421 162 422
rect 162 421 163 422
rect 163 421 164 422
rect 164 421 165 422
rect 165 421 166 422
rect 461 421 462 422
rect 462 421 463 422
rect 463 421 464 422
rect 464 421 465 422
rect 465 421 466 422
rect 466 421 467 422
rect 467 421 468 422
rect 468 421 469 422
rect 469 421 470 422
rect 470 421 471 422
rect 471 421 472 422
rect 104 420 105 421
rect 105 420 106 421
rect 106 420 107 421
rect 107 420 108 421
rect 108 420 109 421
rect 109 420 110 421
rect 110 420 111 421
rect 111 420 112 421
rect 112 420 113 421
rect 113 420 114 421
rect 114 420 115 421
rect 115 420 116 421
rect 116 420 117 421
rect 117 420 118 421
rect 118 420 119 421
rect 119 420 120 421
rect 120 420 121 421
rect 121 420 122 421
rect 122 420 123 421
rect 123 420 124 421
rect 124 420 125 421
rect 125 420 126 421
rect 126 420 127 421
rect 127 420 128 421
rect 128 420 129 421
rect 129 420 130 421
rect 130 420 131 421
rect 131 420 132 421
rect 132 420 133 421
rect 133 420 134 421
rect 134 420 135 421
rect 135 420 136 421
rect 136 420 137 421
rect 137 420 138 421
rect 138 420 139 421
rect 150 420 151 421
rect 151 420 152 421
rect 152 420 153 421
rect 153 420 154 421
rect 154 420 155 421
rect 155 420 156 421
rect 156 420 157 421
rect 157 420 158 421
rect 158 420 159 421
rect 159 420 160 421
rect 160 420 161 421
rect 161 420 162 421
rect 162 420 163 421
rect 163 420 164 421
rect 164 420 165 421
rect 462 420 463 421
rect 463 420 464 421
rect 464 420 465 421
rect 465 420 466 421
rect 466 420 467 421
rect 467 420 468 421
rect 468 420 469 421
rect 469 420 470 421
rect 470 420 471 421
rect 471 420 472 421
rect 472 420 473 421
rect 101 419 102 420
rect 102 419 103 420
rect 103 419 104 420
rect 104 419 105 420
rect 105 419 106 420
rect 106 419 107 420
rect 107 419 108 420
rect 108 419 109 420
rect 109 419 110 420
rect 110 419 111 420
rect 111 419 112 420
rect 112 419 113 420
rect 113 419 114 420
rect 114 419 115 420
rect 115 419 116 420
rect 116 419 117 420
rect 117 419 118 420
rect 118 419 119 420
rect 119 419 120 420
rect 120 419 121 420
rect 121 419 122 420
rect 122 419 123 420
rect 123 419 124 420
rect 124 419 125 420
rect 125 419 126 420
rect 126 419 127 420
rect 127 419 128 420
rect 128 419 129 420
rect 129 419 130 420
rect 130 419 131 420
rect 131 419 132 420
rect 132 419 133 420
rect 133 419 134 420
rect 134 419 135 420
rect 135 419 136 420
rect 136 419 137 420
rect 137 419 138 420
rect 138 419 139 420
rect 139 419 140 420
rect 140 419 141 420
rect 141 419 142 420
rect 150 419 151 420
rect 151 419 152 420
rect 152 419 153 420
rect 153 419 154 420
rect 154 419 155 420
rect 155 419 156 420
rect 156 419 157 420
rect 157 419 158 420
rect 158 419 159 420
rect 159 419 160 420
rect 160 419 161 420
rect 161 419 162 420
rect 162 419 163 420
rect 163 419 164 420
rect 463 419 464 420
rect 464 419 465 420
rect 465 419 466 420
rect 466 419 467 420
rect 467 419 468 420
rect 468 419 469 420
rect 469 419 470 420
rect 470 419 471 420
rect 471 419 472 420
rect 472 419 473 420
rect 473 419 474 420
rect 99 418 100 419
rect 100 418 101 419
rect 101 418 102 419
rect 102 418 103 419
rect 103 418 104 419
rect 104 418 105 419
rect 105 418 106 419
rect 106 418 107 419
rect 107 418 108 419
rect 108 418 109 419
rect 109 418 110 419
rect 110 418 111 419
rect 111 418 112 419
rect 112 418 113 419
rect 113 418 114 419
rect 114 418 115 419
rect 115 418 116 419
rect 116 418 117 419
rect 117 418 118 419
rect 118 418 119 419
rect 119 418 120 419
rect 120 418 121 419
rect 121 418 122 419
rect 122 418 123 419
rect 123 418 124 419
rect 124 418 125 419
rect 125 418 126 419
rect 126 418 127 419
rect 127 418 128 419
rect 128 418 129 419
rect 129 418 130 419
rect 130 418 131 419
rect 131 418 132 419
rect 132 418 133 419
rect 133 418 134 419
rect 134 418 135 419
rect 135 418 136 419
rect 136 418 137 419
rect 137 418 138 419
rect 138 418 139 419
rect 139 418 140 419
rect 140 418 141 419
rect 141 418 142 419
rect 142 418 143 419
rect 143 418 144 419
rect 144 418 145 419
rect 148 418 149 419
rect 149 418 150 419
rect 150 418 151 419
rect 151 418 152 419
rect 152 418 153 419
rect 153 418 154 419
rect 154 418 155 419
rect 155 418 156 419
rect 156 418 157 419
rect 157 418 158 419
rect 158 418 159 419
rect 159 418 160 419
rect 160 418 161 419
rect 161 418 162 419
rect 162 418 163 419
rect 464 418 465 419
rect 465 418 466 419
rect 466 418 467 419
rect 467 418 468 419
rect 468 418 469 419
rect 469 418 470 419
rect 470 418 471 419
rect 471 418 472 419
rect 472 418 473 419
rect 473 418 474 419
rect 474 418 475 419
rect 97 417 98 418
rect 98 417 99 418
rect 99 417 100 418
rect 100 417 101 418
rect 101 417 102 418
rect 102 417 103 418
rect 103 417 104 418
rect 104 417 105 418
rect 105 417 106 418
rect 106 417 107 418
rect 107 417 108 418
rect 108 417 109 418
rect 109 417 110 418
rect 110 417 111 418
rect 111 417 112 418
rect 112 417 113 418
rect 113 417 114 418
rect 114 417 115 418
rect 115 417 116 418
rect 116 417 117 418
rect 117 417 118 418
rect 118 417 119 418
rect 119 417 120 418
rect 120 417 121 418
rect 121 417 122 418
rect 122 417 123 418
rect 123 417 124 418
rect 124 417 125 418
rect 125 417 126 418
rect 126 417 127 418
rect 127 417 128 418
rect 128 417 129 418
rect 129 417 130 418
rect 130 417 131 418
rect 131 417 132 418
rect 132 417 133 418
rect 133 417 134 418
rect 134 417 135 418
rect 135 417 136 418
rect 136 417 137 418
rect 137 417 138 418
rect 138 417 139 418
rect 139 417 140 418
rect 140 417 141 418
rect 141 417 142 418
rect 142 417 143 418
rect 143 417 144 418
rect 144 417 145 418
rect 145 417 146 418
rect 146 417 147 418
rect 147 417 148 418
rect 148 417 149 418
rect 149 417 150 418
rect 150 417 151 418
rect 151 417 152 418
rect 152 417 153 418
rect 153 417 154 418
rect 154 417 155 418
rect 155 417 156 418
rect 156 417 157 418
rect 157 417 158 418
rect 158 417 159 418
rect 159 417 160 418
rect 160 417 161 418
rect 465 417 466 418
rect 466 417 467 418
rect 467 417 468 418
rect 468 417 469 418
rect 469 417 470 418
rect 470 417 471 418
rect 471 417 472 418
rect 472 417 473 418
rect 473 417 474 418
rect 474 417 475 418
rect 475 417 476 418
rect 95 416 96 417
rect 96 416 97 417
rect 97 416 98 417
rect 98 416 99 417
rect 99 416 100 417
rect 100 416 101 417
rect 101 416 102 417
rect 102 416 103 417
rect 103 416 104 417
rect 104 416 105 417
rect 105 416 106 417
rect 106 416 107 417
rect 107 416 108 417
rect 108 416 109 417
rect 109 416 110 417
rect 110 416 111 417
rect 111 416 112 417
rect 112 416 113 417
rect 113 416 114 417
rect 114 416 115 417
rect 115 416 116 417
rect 116 416 117 417
rect 117 416 118 417
rect 118 416 119 417
rect 119 416 120 417
rect 120 416 121 417
rect 121 416 122 417
rect 122 416 123 417
rect 123 416 124 417
rect 124 416 125 417
rect 125 416 126 417
rect 126 416 127 417
rect 127 416 128 417
rect 128 416 129 417
rect 129 416 130 417
rect 130 416 131 417
rect 131 416 132 417
rect 132 416 133 417
rect 133 416 134 417
rect 134 416 135 417
rect 135 416 136 417
rect 136 416 137 417
rect 137 416 138 417
rect 138 416 139 417
rect 139 416 140 417
rect 140 416 141 417
rect 141 416 142 417
rect 142 416 143 417
rect 143 416 144 417
rect 144 416 145 417
rect 145 416 146 417
rect 146 416 147 417
rect 147 416 148 417
rect 148 416 149 417
rect 149 416 150 417
rect 150 416 151 417
rect 151 416 152 417
rect 152 416 153 417
rect 153 416 154 417
rect 154 416 155 417
rect 155 416 156 417
rect 156 416 157 417
rect 157 416 158 417
rect 158 416 159 417
rect 159 416 160 417
rect 466 416 467 417
rect 467 416 468 417
rect 468 416 469 417
rect 469 416 470 417
rect 470 416 471 417
rect 471 416 472 417
rect 472 416 473 417
rect 473 416 474 417
rect 474 416 475 417
rect 475 416 476 417
rect 476 416 477 417
rect 94 415 95 416
rect 95 415 96 416
rect 96 415 97 416
rect 97 415 98 416
rect 98 415 99 416
rect 99 415 100 416
rect 100 415 101 416
rect 101 415 102 416
rect 102 415 103 416
rect 103 415 104 416
rect 104 415 105 416
rect 105 415 106 416
rect 106 415 107 416
rect 107 415 108 416
rect 108 415 109 416
rect 109 415 110 416
rect 110 415 111 416
rect 111 415 112 416
rect 112 415 113 416
rect 113 415 114 416
rect 114 415 115 416
rect 115 415 116 416
rect 116 415 117 416
rect 117 415 118 416
rect 118 415 119 416
rect 119 415 120 416
rect 120 415 121 416
rect 121 415 122 416
rect 122 415 123 416
rect 123 415 124 416
rect 124 415 125 416
rect 125 415 126 416
rect 126 415 127 416
rect 127 415 128 416
rect 128 415 129 416
rect 129 415 130 416
rect 130 415 131 416
rect 131 415 132 416
rect 132 415 133 416
rect 133 415 134 416
rect 134 415 135 416
rect 135 415 136 416
rect 136 415 137 416
rect 137 415 138 416
rect 138 415 139 416
rect 139 415 140 416
rect 140 415 141 416
rect 141 415 142 416
rect 142 415 143 416
rect 143 415 144 416
rect 144 415 145 416
rect 145 415 146 416
rect 146 415 147 416
rect 147 415 148 416
rect 148 415 149 416
rect 149 415 150 416
rect 150 415 151 416
rect 151 415 152 416
rect 152 415 153 416
rect 153 415 154 416
rect 154 415 155 416
rect 155 415 156 416
rect 156 415 157 416
rect 157 415 158 416
rect 158 415 159 416
rect 467 415 468 416
rect 468 415 469 416
rect 469 415 470 416
rect 470 415 471 416
rect 471 415 472 416
rect 472 415 473 416
rect 473 415 474 416
rect 474 415 475 416
rect 475 415 476 416
rect 476 415 477 416
rect 477 415 478 416
rect 92 414 93 415
rect 93 414 94 415
rect 94 414 95 415
rect 95 414 96 415
rect 96 414 97 415
rect 97 414 98 415
rect 98 414 99 415
rect 99 414 100 415
rect 100 414 101 415
rect 101 414 102 415
rect 102 414 103 415
rect 103 414 104 415
rect 104 414 105 415
rect 105 414 106 415
rect 106 414 107 415
rect 107 414 108 415
rect 108 414 109 415
rect 109 414 110 415
rect 110 414 111 415
rect 111 414 112 415
rect 112 414 113 415
rect 113 414 114 415
rect 114 414 115 415
rect 115 414 116 415
rect 125 414 126 415
rect 126 414 127 415
rect 127 414 128 415
rect 128 414 129 415
rect 129 414 130 415
rect 130 414 131 415
rect 131 414 132 415
rect 132 414 133 415
rect 133 414 134 415
rect 134 414 135 415
rect 135 414 136 415
rect 136 414 137 415
rect 137 414 138 415
rect 138 414 139 415
rect 139 414 140 415
rect 140 414 141 415
rect 141 414 142 415
rect 142 414 143 415
rect 143 414 144 415
rect 144 414 145 415
rect 145 414 146 415
rect 146 414 147 415
rect 147 414 148 415
rect 148 414 149 415
rect 149 414 150 415
rect 150 414 151 415
rect 151 414 152 415
rect 152 414 153 415
rect 153 414 154 415
rect 154 414 155 415
rect 155 414 156 415
rect 156 414 157 415
rect 157 414 158 415
rect 468 414 469 415
rect 469 414 470 415
rect 470 414 471 415
rect 471 414 472 415
rect 472 414 473 415
rect 473 414 474 415
rect 474 414 475 415
rect 475 414 476 415
rect 476 414 477 415
rect 477 414 478 415
rect 478 414 479 415
rect 91 413 92 414
rect 92 413 93 414
rect 93 413 94 414
rect 94 413 95 414
rect 95 413 96 414
rect 96 413 97 414
rect 97 413 98 414
rect 98 413 99 414
rect 99 413 100 414
rect 100 413 101 414
rect 101 413 102 414
rect 102 413 103 414
rect 103 413 104 414
rect 104 413 105 414
rect 105 413 106 414
rect 106 413 107 414
rect 107 413 108 414
rect 108 413 109 414
rect 109 413 110 414
rect 110 413 111 414
rect 132 413 133 414
rect 133 413 134 414
rect 134 413 135 414
rect 135 413 136 414
rect 136 413 137 414
rect 137 413 138 414
rect 138 413 139 414
rect 139 413 140 414
rect 140 413 141 414
rect 141 413 142 414
rect 142 413 143 414
rect 143 413 144 414
rect 144 413 145 414
rect 145 413 146 414
rect 146 413 147 414
rect 147 413 148 414
rect 148 413 149 414
rect 149 413 150 414
rect 150 413 151 414
rect 151 413 152 414
rect 152 413 153 414
rect 153 413 154 414
rect 154 413 155 414
rect 155 413 156 414
rect 468 413 469 414
rect 469 413 470 414
rect 470 413 471 414
rect 471 413 472 414
rect 472 413 473 414
rect 473 413 474 414
rect 474 413 475 414
rect 475 413 476 414
rect 476 413 477 414
rect 477 413 478 414
rect 478 413 479 414
rect 479 413 480 414
rect 90 412 91 413
rect 91 412 92 413
rect 92 412 93 413
rect 93 412 94 413
rect 94 412 95 413
rect 95 412 96 413
rect 96 412 97 413
rect 97 412 98 413
rect 98 412 99 413
rect 99 412 100 413
rect 100 412 101 413
rect 101 412 102 413
rect 102 412 103 413
rect 103 412 104 413
rect 104 412 105 413
rect 105 412 106 413
rect 106 412 107 413
rect 107 412 108 413
rect 136 412 137 413
rect 137 412 138 413
rect 138 412 139 413
rect 139 412 140 413
rect 140 412 141 413
rect 141 412 142 413
rect 142 412 143 413
rect 143 412 144 413
rect 144 412 145 413
rect 145 412 146 413
rect 146 412 147 413
rect 147 412 148 413
rect 148 412 149 413
rect 149 412 150 413
rect 150 412 151 413
rect 151 412 152 413
rect 152 412 153 413
rect 153 412 154 413
rect 154 412 155 413
rect 469 412 470 413
rect 470 412 471 413
rect 471 412 472 413
rect 472 412 473 413
rect 473 412 474 413
rect 474 412 475 413
rect 475 412 476 413
rect 476 412 477 413
rect 477 412 478 413
rect 478 412 479 413
rect 479 412 480 413
rect 480 412 481 413
rect 88 411 89 412
rect 89 411 90 412
rect 90 411 91 412
rect 91 411 92 412
rect 92 411 93 412
rect 93 411 94 412
rect 94 411 95 412
rect 95 411 96 412
rect 96 411 97 412
rect 97 411 98 412
rect 98 411 99 412
rect 99 411 100 412
rect 100 411 101 412
rect 101 411 102 412
rect 102 411 103 412
rect 103 411 104 412
rect 104 411 105 412
rect 139 411 140 412
rect 140 411 141 412
rect 141 411 142 412
rect 142 411 143 412
rect 143 411 144 412
rect 144 411 145 412
rect 145 411 146 412
rect 146 411 147 412
rect 147 411 148 412
rect 148 411 149 412
rect 149 411 150 412
rect 150 411 151 412
rect 151 411 152 412
rect 152 411 153 412
rect 153 411 154 412
rect 470 411 471 412
rect 471 411 472 412
rect 472 411 473 412
rect 473 411 474 412
rect 474 411 475 412
rect 475 411 476 412
rect 476 411 477 412
rect 477 411 478 412
rect 478 411 479 412
rect 479 411 480 412
rect 480 411 481 412
rect 481 411 482 412
rect 87 410 88 411
rect 88 410 89 411
rect 89 410 90 411
rect 90 410 91 411
rect 91 410 92 411
rect 92 410 93 411
rect 93 410 94 411
rect 94 410 95 411
rect 95 410 96 411
rect 96 410 97 411
rect 97 410 98 411
rect 98 410 99 411
rect 99 410 100 411
rect 100 410 101 411
rect 101 410 102 411
rect 102 410 103 411
rect 141 410 142 411
rect 142 410 143 411
rect 143 410 144 411
rect 144 410 145 411
rect 145 410 146 411
rect 146 410 147 411
rect 147 410 148 411
rect 148 410 149 411
rect 149 410 150 411
rect 150 410 151 411
rect 151 410 152 411
rect 233 410 234 411
rect 234 410 235 411
rect 235 410 236 411
rect 236 410 237 411
rect 237 410 238 411
rect 238 410 239 411
rect 239 410 240 411
rect 240 410 241 411
rect 241 410 242 411
rect 242 410 243 411
rect 243 410 244 411
rect 244 410 245 411
rect 245 410 246 411
rect 246 410 247 411
rect 247 410 248 411
rect 248 410 249 411
rect 471 410 472 411
rect 472 410 473 411
rect 473 410 474 411
rect 474 410 475 411
rect 475 410 476 411
rect 476 410 477 411
rect 477 410 478 411
rect 478 410 479 411
rect 479 410 480 411
rect 480 410 481 411
rect 481 410 482 411
rect 482 410 483 411
rect 86 409 87 410
rect 87 409 88 410
rect 88 409 89 410
rect 89 409 90 410
rect 90 409 91 410
rect 91 409 92 410
rect 92 409 93 410
rect 93 409 94 410
rect 94 409 95 410
rect 95 409 96 410
rect 96 409 97 410
rect 97 409 98 410
rect 98 409 99 410
rect 99 409 100 410
rect 100 409 101 410
rect 140 409 141 410
rect 141 409 142 410
rect 142 409 143 410
rect 143 409 144 410
rect 144 409 145 410
rect 145 409 146 410
rect 146 409 147 410
rect 147 409 148 410
rect 148 409 149 410
rect 149 409 150 410
rect 150 409 151 410
rect 228 409 229 410
rect 229 409 230 410
rect 230 409 231 410
rect 231 409 232 410
rect 232 409 233 410
rect 233 409 234 410
rect 234 409 235 410
rect 235 409 236 410
rect 236 409 237 410
rect 237 409 238 410
rect 238 409 239 410
rect 239 409 240 410
rect 240 409 241 410
rect 241 409 242 410
rect 242 409 243 410
rect 243 409 244 410
rect 244 409 245 410
rect 245 409 246 410
rect 246 409 247 410
rect 247 409 248 410
rect 248 409 249 410
rect 249 409 250 410
rect 250 409 251 410
rect 251 409 252 410
rect 252 409 253 410
rect 253 409 254 410
rect 472 409 473 410
rect 473 409 474 410
rect 474 409 475 410
rect 475 409 476 410
rect 476 409 477 410
rect 477 409 478 410
rect 478 409 479 410
rect 479 409 480 410
rect 480 409 481 410
rect 481 409 482 410
rect 482 409 483 410
rect 85 408 86 409
rect 86 408 87 409
rect 87 408 88 409
rect 88 408 89 409
rect 89 408 90 409
rect 90 408 91 409
rect 91 408 92 409
rect 92 408 93 409
rect 93 408 94 409
rect 94 408 95 409
rect 95 408 96 409
rect 96 408 97 409
rect 97 408 98 409
rect 98 408 99 409
rect 139 408 140 409
rect 140 408 141 409
rect 141 408 142 409
rect 142 408 143 409
rect 143 408 144 409
rect 144 408 145 409
rect 145 408 146 409
rect 146 408 147 409
rect 147 408 148 409
rect 148 408 149 409
rect 149 408 150 409
rect 224 408 225 409
rect 225 408 226 409
rect 226 408 227 409
rect 227 408 228 409
rect 228 408 229 409
rect 229 408 230 409
rect 230 408 231 409
rect 231 408 232 409
rect 232 408 233 409
rect 233 408 234 409
rect 234 408 235 409
rect 235 408 236 409
rect 236 408 237 409
rect 237 408 238 409
rect 238 408 239 409
rect 239 408 240 409
rect 240 408 241 409
rect 241 408 242 409
rect 242 408 243 409
rect 243 408 244 409
rect 244 408 245 409
rect 245 408 246 409
rect 246 408 247 409
rect 247 408 248 409
rect 248 408 249 409
rect 249 408 250 409
rect 250 408 251 409
rect 251 408 252 409
rect 252 408 253 409
rect 253 408 254 409
rect 254 408 255 409
rect 255 408 256 409
rect 256 408 257 409
rect 473 408 474 409
rect 474 408 475 409
rect 475 408 476 409
rect 476 408 477 409
rect 477 408 478 409
rect 478 408 479 409
rect 479 408 480 409
rect 480 408 481 409
rect 481 408 482 409
rect 482 408 483 409
rect 483 408 484 409
rect 84 407 85 408
rect 85 407 86 408
rect 86 407 87 408
rect 87 407 88 408
rect 88 407 89 408
rect 89 407 90 408
rect 90 407 91 408
rect 91 407 92 408
rect 92 407 93 408
rect 93 407 94 408
rect 94 407 95 408
rect 95 407 96 408
rect 96 407 97 408
rect 97 407 98 408
rect 138 407 139 408
rect 139 407 140 408
rect 140 407 141 408
rect 141 407 142 408
rect 142 407 143 408
rect 143 407 144 408
rect 144 407 145 408
rect 145 407 146 408
rect 146 407 147 408
rect 147 407 148 408
rect 220 407 221 408
rect 221 407 222 408
rect 222 407 223 408
rect 223 407 224 408
rect 224 407 225 408
rect 225 407 226 408
rect 226 407 227 408
rect 227 407 228 408
rect 228 407 229 408
rect 229 407 230 408
rect 230 407 231 408
rect 231 407 232 408
rect 232 407 233 408
rect 233 407 234 408
rect 234 407 235 408
rect 235 407 236 408
rect 236 407 237 408
rect 237 407 238 408
rect 238 407 239 408
rect 239 407 240 408
rect 240 407 241 408
rect 241 407 242 408
rect 242 407 243 408
rect 243 407 244 408
rect 244 407 245 408
rect 245 407 246 408
rect 246 407 247 408
rect 247 407 248 408
rect 248 407 249 408
rect 249 407 250 408
rect 250 407 251 408
rect 251 407 252 408
rect 252 407 253 408
rect 253 407 254 408
rect 254 407 255 408
rect 255 407 256 408
rect 256 407 257 408
rect 257 407 258 408
rect 258 407 259 408
rect 259 407 260 408
rect 474 407 475 408
rect 475 407 476 408
rect 476 407 477 408
rect 477 407 478 408
rect 478 407 479 408
rect 479 407 480 408
rect 480 407 481 408
rect 481 407 482 408
rect 482 407 483 408
rect 483 407 484 408
rect 484 407 485 408
rect 83 406 84 407
rect 84 406 85 407
rect 85 406 86 407
rect 86 406 87 407
rect 87 406 88 407
rect 88 406 89 407
rect 89 406 90 407
rect 90 406 91 407
rect 91 406 92 407
rect 92 406 93 407
rect 93 406 94 407
rect 94 406 95 407
rect 95 406 96 407
rect 137 406 138 407
rect 138 406 139 407
rect 139 406 140 407
rect 140 406 141 407
rect 141 406 142 407
rect 142 406 143 407
rect 143 406 144 407
rect 144 406 145 407
rect 145 406 146 407
rect 146 406 147 407
rect 218 406 219 407
rect 219 406 220 407
rect 220 406 221 407
rect 221 406 222 407
rect 222 406 223 407
rect 223 406 224 407
rect 224 406 225 407
rect 225 406 226 407
rect 226 406 227 407
rect 227 406 228 407
rect 228 406 229 407
rect 229 406 230 407
rect 230 406 231 407
rect 231 406 232 407
rect 232 406 233 407
rect 233 406 234 407
rect 234 406 235 407
rect 235 406 236 407
rect 236 406 237 407
rect 237 406 238 407
rect 238 406 239 407
rect 239 406 240 407
rect 240 406 241 407
rect 241 406 242 407
rect 242 406 243 407
rect 243 406 244 407
rect 244 406 245 407
rect 245 406 246 407
rect 246 406 247 407
rect 247 406 248 407
rect 248 406 249 407
rect 249 406 250 407
rect 250 406 251 407
rect 251 406 252 407
rect 252 406 253 407
rect 253 406 254 407
rect 254 406 255 407
rect 255 406 256 407
rect 256 406 257 407
rect 257 406 258 407
rect 258 406 259 407
rect 259 406 260 407
rect 260 406 261 407
rect 261 406 262 407
rect 475 406 476 407
rect 476 406 477 407
rect 477 406 478 407
rect 478 406 479 407
rect 479 406 480 407
rect 480 406 481 407
rect 481 406 482 407
rect 482 406 483 407
rect 483 406 484 407
rect 484 406 485 407
rect 82 405 83 406
rect 83 405 84 406
rect 84 405 85 406
rect 85 405 86 406
rect 86 405 87 406
rect 87 405 88 406
rect 88 405 89 406
rect 89 405 90 406
rect 90 405 91 406
rect 91 405 92 406
rect 92 405 93 406
rect 93 405 94 406
rect 94 405 95 406
rect 135 405 136 406
rect 136 405 137 406
rect 137 405 138 406
rect 138 405 139 406
rect 139 405 140 406
rect 140 405 141 406
rect 141 405 142 406
rect 142 405 143 406
rect 143 405 144 406
rect 144 405 145 406
rect 216 405 217 406
rect 217 405 218 406
rect 218 405 219 406
rect 219 405 220 406
rect 220 405 221 406
rect 221 405 222 406
rect 222 405 223 406
rect 223 405 224 406
rect 224 405 225 406
rect 225 405 226 406
rect 226 405 227 406
rect 227 405 228 406
rect 228 405 229 406
rect 229 405 230 406
rect 230 405 231 406
rect 231 405 232 406
rect 232 405 233 406
rect 233 405 234 406
rect 234 405 235 406
rect 235 405 236 406
rect 236 405 237 406
rect 237 405 238 406
rect 238 405 239 406
rect 239 405 240 406
rect 240 405 241 406
rect 241 405 242 406
rect 242 405 243 406
rect 243 405 244 406
rect 244 405 245 406
rect 245 405 246 406
rect 246 405 247 406
rect 247 405 248 406
rect 248 405 249 406
rect 249 405 250 406
rect 250 405 251 406
rect 251 405 252 406
rect 252 405 253 406
rect 253 405 254 406
rect 254 405 255 406
rect 255 405 256 406
rect 256 405 257 406
rect 257 405 258 406
rect 258 405 259 406
rect 259 405 260 406
rect 260 405 261 406
rect 261 405 262 406
rect 262 405 263 406
rect 263 405 264 406
rect 476 405 477 406
rect 477 405 478 406
rect 478 405 479 406
rect 479 405 480 406
rect 480 405 481 406
rect 481 405 482 406
rect 482 405 483 406
rect 483 405 484 406
rect 484 405 485 406
rect 485 405 486 406
rect 81 404 82 405
rect 82 404 83 405
rect 83 404 84 405
rect 84 404 85 405
rect 85 404 86 405
rect 86 404 87 405
rect 87 404 88 405
rect 88 404 89 405
rect 89 404 90 405
rect 90 404 91 405
rect 91 404 92 405
rect 92 404 93 405
rect 93 404 94 405
rect 134 404 135 405
rect 135 404 136 405
rect 136 404 137 405
rect 137 404 138 405
rect 138 404 139 405
rect 139 404 140 405
rect 140 404 141 405
rect 141 404 142 405
rect 142 404 143 405
rect 214 404 215 405
rect 215 404 216 405
rect 216 404 217 405
rect 217 404 218 405
rect 218 404 219 405
rect 219 404 220 405
rect 220 404 221 405
rect 221 404 222 405
rect 222 404 223 405
rect 223 404 224 405
rect 224 404 225 405
rect 225 404 226 405
rect 226 404 227 405
rect 227 404 228 405
rect 228 404 229 405
rect 229 404 230 405
rect 230 404 231 405
rect 231 404 232 405
rect 232 404 233 405
rect 233 404 234 405
rect 234 404 235 405
rect 235 404 236 405
rect 236 404 237 405
rect 237 404 238 405
rect 238 404 239 405
rect 239 404 240 405
rect 240 404 241 405
rect 241 404 242 405
rect 242 404 243 405
rect 243 404 244 405
rect 244 404 245 405
rect 245 404 246 405
rect 246 404 247 405
rect 247 404 248 405
rect 248 404 249 405
rect 249 404 250 405
rect 250 404 251 405
rect 251 404 252 405
rect 252 404 253 405
rect 253 404 254 405
rect 254 404 255 405
rect 255 404 256 405
rect 256 404 257 405
rect 257 404 258 405
rect 258 404 259 405
rect 259 404 260 405
rect 260 404 261 405
rect 261 404 262 405
rect 262 404 263 405
rect 263 404 264 405
rect 264 404 265 405
rect 477 404 478 405
rect 478 404 479 405
rect 479 404 480 405
rect 480 404 481 405
rect 481 404 482 405
rect 482 404 483 405
rect 483 404 484 405
rect 484 404 485 405
rect 485 404 486 405
rect 486 404 487 405
rect 80 403 81 404
rect 81 403 82 404
rect 82 403 83 404
rect 83 403 84 404
rect 84 403 85 404
rect 85 403 86 404
rect 86 403 87 404
rect 87 403 88 404
rect 88 403 89 404
rect 89 403 90 404
rect 90 403 91 404
rect 91 403 92 404
rect 92 403 93 404
rect 132 403 133 404
rect 133 403 134 404
rect 134 403 135 404
rect 135 403 136 404
rect 136 403 137 404
rect 137 403 138 404
rect 138 403 139 404
rect 139 403 140 404
rect 140 403 141 404
rect 141 403 142 404
rect 212 403 213 404
rect 213 403 214 404
rect 214 403 215 404
rect 215 403 216 404
rect 216 403 217 404
rect 217 403 218 404
rect 218 403 219 404
rect 219 403 220 404
rect 220 403 221 404
rect 221 403 222 404
rect 222 403 223 404
rect 223 403 224 404
rect 224 403 225 404
rect 225 403 226 404
rect 226 403 227 404
rect 227 403 228 404
rect 228 403 229 404
rect 229 403 230 404
rect 230 403 231 404
rect 231 403 232 404
rect 232 403 233 404
rect 233 403 234 404
rect 234 403 235 404
rect 235 403 236 404
rect 236 403 237 404
rect 237 403 238 404
rect 238 403 239 404
rect 239 403 240 404
rect 240 403 241 404
rect 241 403 242 404
rect 242 403 243 404
rect 243 403 244 404
rect 244 403 245 404
rect 245 403 246 404
rect 246 403 247 404
rect 247 403 248 404
rect 248 403 249 404
rect 249 403 250 404
rect 250 403 251 404
rect 251 403 252 404
rect 252 403 253 404
rect 253 403 254 404
rect 254 403 255 404
rect 255 403 256 404
rect 256 403 257 404
rect 257 403 258 404
rect 258 403 259 404
rect 259 403 260 404
rect 260 403 261 404
rect 261 403 262 404
rect 262 403 263 404
rect 263 403 264 404
rect 264 403 265 404
rect 265 403 266 404
rect 266 403 267 404
rect 477 403 478 404
rect 478 403 479 404
rect 479 403 480 404
rect 480 403 481 404
rect 481 403 482 404
rect 482 403 483 404
rect 483 403 484 404
rect 484 403 485 404
rect 485 403 486 404
rect 486 403 487 404
rect 79 402 80 403
rect 80 402 81 403
rect 81 402 82 403
rect 82 402 83 403
rect 83 402 84 403
rect 84 402 85 403
rect 85 402 86 403
rect 86 402 87 403
rect 87 402 88 403
rect 88 402 89 403
rect 89 402 90 403
rect 90 402 91 403
rect 91 402 92 403
rect 131 402 132 403
rect 132 402 133 403
rect 133 402 134 403
rect 134 402 135 403
rect 135 402 136 403
rect 136 402 137 403
rect 137 402 138 403
rect 138 402 139 403
rect 139 402 140 403
rect 210 402 211 403
rect 211 402 212 403
rect 212 402 213 403
rect 213 402 214 403
rect 214 402 215 403
rect 215 402 216 403
rect 216 402 217 403
rect 217 402 218 403
rect 218 402 219 403
rect 219 402 220 403
rect 220 402 221 403
rect 221 402 222 403
rect 222 402 223 403
rect 223 402 224 403
rect 224 402 225 403
rect 225 402 226 403
rect 226 402 227 403
rect 227 402 228 403
rect 228 402 229 403
rect 229 402 230 403
rect 230 402 231 403
rect 231 402 232 403
rect 232 402 233 403
rect 233 402 234 403
rect 234 402 235 403
rect 235 402 236 403
rect 236 402 237 403
rect 237 402 238 403
rect 238 402 239 403
rect 239 402 240 403
rect 240 402 241 403
rect 241 402 242 403
rect 242 402 243 403
rect 243 402 244 403
rect 244 402 245 403
rect 245 402 246 403
rect 246 402 247 403
rect 247 402 248 403
rect 248 402 249 403
rect 249 402 250 403
rect 250 402 251 403
rect 251 402 252 403
rect 252 402 253 403
rect 253 402 254 403
rect 254 402 255 403
rect 255 402 256 403
rect 256 402 257 403
rect 257 402 258 403
rect 258 402 259 403
rect 259 402 260 403
rect 260 402 261 403
rect 261 402 262 403
rect 262 402 263 403
rect 263 402 264 403
rect 264 402 265 403
rect 265 402 266 403
rect 266 402 267 403
rect 267 402 268 403
rect 478 402 479 403
rect 479 402 480 403
rect 480 402 481 403
rect 481 402 482 403
rect 482 402 483 403
rect 483 402 484 403
rect 484 402 485 403
rect 485 402 486 403
rect 486 402 487 403
rect 487 402 488 403
rect 79 401 80 402
rect 80 401 81 402
rect 81 401 82 402
rect 82 401 83 402
rect 83 401 84 402
rect 84 401 85 402
rect 85 401 86 402
rect 86 401 87 402
rect 87 401 88 402
rect 88 401 89 402
rect 89 401 90 402
rect 90 401 91 402
rect 129 401 130 402
rect 130 401 131 402
rect 131 401 132 402
rect 132 401 133 402
rect 133 401 134 402
rect 134 401 135 402
rect 135 401 136 402
rect 136 401 137 402
rect 137 401 138 402
rect 209 401 210 402
rect 210 401 211 402
rect 211 401 212 402
rect 212 401 213 402
rect 213 401 214 402
rect 214 401 215 402
rect 215 401 216 402
rect 216 401 217 402
rect 217 401 218 402
rect 218 401 219 402
rect 219 401 220 402
rect 220 401 221 402
rect 221 401 222 402
rect 222 401 223 402
rect 223 401 224 402
rect 224 401 225 402
rect 225 401 226 402
rect 226 401 227 402
rect 227 401 228 402
rect 228 401 229 402
rect 229 401 230 402
rect 230 401 231 402
rect 231 401 232 402
rect 232 401 233 402
rect 233 401 234 402
rect 234 401 235 402
rect 235 401 236 402
rect 236 401 237 402
rect 237 401 238 402
rect 238 401 239 402
rect 239 401 240 402
rect 240 401 241 402
rect 241 401 242 402
rect 242 401 243 402
rect 243 401 244 402
rect 244 401 245 402
rect 245 401 246 402
rect 246 401 247 402
rect 247 401 248 402
rect 248 401 249 402
rect 249 401 250 402
rect 250 401 251 402
rect 251 401 252 402
rect 252 401 253 402
rect 253 401 254 402
rect 254 401 255 402
rect 255 401 256 402
rect 256 401 257 402
rect 257 401 258 402
rect 258 401 259 402
rect 259 401 260 402
rect 260 401 261 402
rect 261 401 262 402
rect 262 401 263 402
rect 263 401 264 402
rect 264 401 265 402
rect 265 401 266 402
rect 266 401 267 402
rect 267 401 268 402
rect 268 401 269 402
rect 269 401 270 402
rect 479 401 480 402
rect 480 401 481 402
rect 481 401 482 402
rect 482 401 483 402
rect 483 401 484 402
rect 484 401 485 402
rect 485 401 486 402
rect 486 401 487 402
rect 487 401 488 402
rect 78 400 79 401
rect 79 400 80 401
rect 80 400 81 401
rect 81 400 82 401
rect 82 400 83 401
rect 83 400 84 401
rect 84 400 85 401
rect 85 400 86 401
rect 86 400 87 401
rect 87 400 88 401
rect 88 400 89 401
rect 89 400 90 401
rect 127 400 128 401
rect 128 400 129 401
rect 129 400 130 401
rect 130 400 131 401
rect 131 400 132 401
rect 132 400 133 401
rect 133 400 134 401
rect 134 400 135 401
rect 135 400 136 401
rect 207 400 208 401
rect 208 400 209 401
rect 209 400 210 401
rect 210 400 211 401
rect 211 400 212 401
rect 212 400 213 401
rect 213 400 214 401
rect 214 400 215 401
rect 215 400 216 401
rect 216 400 217 401
rect 217 400 218 401
rect 218 400 219 401
rect 219 400 220 401
rect 220 400 221 401
rect 221 400 222 401
rect 222 400 223 401
rect 223 400 224 401
rect 224 400 225 401
rect 225 400 226 401
rect 226 400 227 401
rect 227 400 228 401
rect 228 400 229 401
rect 229 400 230 401
rect 230 400 231 401
rect 231 400 232 401
rect 232 400 233 401
rect 233 400 234 401
rect 234 400 235 401
rect 235 400 236 401
rect 236 400 237 401
rect 237 400 238 401
rect 238 400 239 401
rect 239 400 240 401
rect 240 400 241 401
rect 241 400 242 401
rect 242 400 243 401
rect 243 400 244 401
rect 244 400 245 401
rect 245 400 246 401
rect 246 400 247 401
rect 247 400 248 401
rect 248 400 249 401
rect 249 400 250 401
rect 250 400 251 401
rect 251 400 252 401
rect 252 400 253 401
rect 253 400 254 401
rect 254 400 255 401
rect 255 400 256 401
rect 256 400 257 401
rect 257 400 258 401
rect 258 400 259 401
rect 259 400 260 401
rect 260 400 261 401
rect 261 400 262 401
rect 262 400 263 401
rect 263 400 264 401
rect 264 400 265 401
rect 265 400 266 401
rect 266 400 267 401
rect 267 400 268 401
rect 268 400 269 401
rect 269 400 270 401
rect 270 400 271 401
rect 479 400 480 401
rect 480 400 481 401
rect 481 400 482 401
rect 482 400 483 401
rect 483 400 484 401
rect 484 400 485 401
rect 485 400 486 401
rect 486 400 487 401
rect 487 400 488 401
rect 488 400 489 401
rect 77 399 78 400
rect 78 399 79 400
rect 79 399 80 400
rect 80 399 81 400
rect 81 399 82 400
rect 82 399 83 400
rect 83 399 84 400
rect 84 399 85 400
rect 85 399 86 400
rect 86 399 87 400
rect 87 399 88 400
rect 88 399 89 400
rect 126 399 127 400
rect 127 399 128 400
rect 128 399 129 400
rect 129 399 130 400
rect 130 399 131 400
rect 131 399 132 400
rect 132 399 133 400
rect 133 399 134 400
rect 206 399 207 400
rect 207 399 208 400
rect 208 399 209 400
rect 209 399 210 400
rect 210 399 211 400
rect 211 399 212 400
rect 212 399 213 400
rect 213 399 214 400
rect 214 399 215 400
rect 215 399 216 400
rect 216 399 217 400
rect 217 399 218 400
rect 218 399 219 400
rect 219 399 220 400
rect 220 399 221 400
rect 221 399 222 400
rect 222 399 223 400
rect 223 399 224 400
rect 224 399 225 400
rect 225 399 226 400
rect 226 399 227 400
rect 227 399 228 400
rect 228 399 229 400
rect 229 399 230 400
rect 230 399 231 400
rect 231 399 232 400
rect 232 399 233 400
rect 233 399 234 400
rect 234 399 235 400
rect 235 399 236 400
rect 236 399 237 400
rect 237 399 238 400
rect 238 399 239 400
rect 239 399 240 400
rect 240 399 241 400
rect 241 399 242 400
rect 242 399 243 400
rect 243 399 244 400
rect 244 399 245 400
rect 245 399 246 400
rect 246 399 247 400
rect 247 399 248 400
rect 248 399 249 400
rect 249 399 250 400
rect 250 399 251 400
rect 251 399 252 400
rect 252 399 253 400
rect 253 399 254 400
rect 254 399 255 400
rect 255 399 256 400
rect 256 399 257 400
rect 257 399 258 400
rect 258 399 259 400
rect 259 399 260 400
rect 260 399 261 400
rect 261 399 262 400
rect 262 399 263 400
rect 263 399 264 400
rect 264 399 265 400
rect 265 399 266 400
rect 266 399 267 400
rect 267 399 268 400
rect 268 399 269 400
rect 269 399 270 400
rect 270 399 271 400
rect 271 399 272 400
rect 480 399 481 400
rect 481 399 482 400
rect 482 399 483 400
rect 483 399 484 400
rect 484 399 485 400
rect 485 399 486 400
rect 486 399 487 400
rect 487 399 488 400
rect 488 399 489 400
rect 76 398 77 399
rect 77 398 78 399
rect 78 398 79 399
rect 79 398 80 399
rect 80 398 81 399
rect 81 398 82 399
rect 82 398 83 399
rect 83 398 84 399
rect 84 398 85 399
rect 85 398 86 399
rect 86 398 87 399
rect 87 398 88 399
rect 124 398 125 399
rect 125 398 126 399
rect 126 398 127 399
rect 127 398 128 399
rect 128 398 129 399
rect 129 398 130 399
rect 130 398 131 399
rect 131 398 132 399
rect 205 398 206 399
rect 206 398 207 399
rect 207 398 208 399
rect 208 398 209 399
rect 209 398 210 399
rect 210 398 211 399
rect 211 398 212 399
rect 212 398 213 399
rect 213 398 214 399
rect 214 398 215 399
rect 215 398 216 399
rect 216 398 217 399
rect 217 398 218 399
rect 218 398 219 399
rect 219 398 220 399
rect 220 398 221 399
rect 221 398 222 399
rect 222 398 223 399
rect 223 398 224 399
rect 224 398 225 399
rect 225 398 226 399
rect 226 398 227 399
rect 227 398 228 399
rect 228 398 229 399
rect 229 398 230 399
rect 230 398 231 399
rect 231 398 232 399
rect 232 398 233 399
rect 233 398 234 399
rect 234 398 235 399
rect 235 398 236 399
rect 236 398 237 399
rect 237 398 238 399
rect 238 398 239 399
rect 239 398 240 399
rect 240 398 241 399
rect 241 398 242 399
rect 242 398 243 399
rect 243 398 244 399
rect 244 398 245 399
rect 245 398 246 399
rect 246 398 247 399
rect 247 398 248 399
rect 248 398 249 399
rect 249 398 250 399
rect 250 398 251 399
rect 251 398 252 399
rect 252 398 253 399
rect 253 398 254 399
rect 254 398 255 399
rect 255 398 256 399
rect 256 398 257 399
rect 257 398 258 399
rect 258 398 259 399
rect 259 398 260 399
rect 260 398 261 399
rect 261 398 262 399
rect 262 398 263 399
rect 263 398 264 399
rect 264 398 265 399
rect 265 398 266 399
rect 266 398 267 399
rect 267 398 268 399
rect 268 398 269 399
rect 269 398 270 399
rect 270 398 271 399
rect 271 398 272 399
rect 272 398 273 399
rect 273 398 274 399
rect 480 398 481 399
rect 481 398 482 399
rect 482 398 483 399
rect 483 398 484 399
rect 484 398 485 399
rect 485 398 486 399
rect 486 398 487 399
rect 487 398 488 399
rect 488 398 489 399
rect 489 398 490 399
rect 76 397 77 398
rect 77 397 78 398
rect 78 397 79 398
rect 79 397 80 398
rect 80 397 81 398
rect 81 397 82 398
rect 82 397 83 398
rect 83 397 84 398
rect 84 397 85 398
rect 85 397 86 398
rect 86 397 87 398
rect 121 397 122 398
rect 122 397 123 398
rect 123 397 124 398
rect 124 397 125 398
rect 125 397 126 398
rect 126 397 127 398
rect 127 397 128 398
rect 128 397 129 398
rect 129 397 130 398
rect 204 397 205 398
rect 205 397 206 398
rect 206 397 207 398
rect 207 397 208 398
rect 208 397 209 398
rect 209 397 210 398
rect 210 397 211 398
rect 211 397 212 398
rect 212 397 213 398
rect 213 397 214 398
rect 214 397 215 398
rect 215 397 216 398
rect 216 397 217 398
rect 230 397 231 398
rect 231 397 232 398
rect 232 397 233 398
rect 233 397 234 398
rect 234 397 235 398
rect 235 397 236 398
rect 236 397 237 398
rect 237 397 238 398
rect 238 397 239 398
rect 239 397 240 398
rect 240 397 241 398
rect 241 397 242 398
rect 242 397 243 398
rect 243 397 244 398
rect 244 397 245 398
rect 245 397 246 398
rect 246 397 247 398
rect 247 397 248 398
rect 248 397 249 398
rect 249 397 250 398
rect 250 397 251 398
rect 251 397 252 398
rect 252 397 253 398
rect 253 397 254 398
rect 254 397 255 398
rect 255 397 256 398
rect 256 397 257 398
rect 257 397 258 398
rect 258 397 259 398
rect 259 397 260 398
rect 260 397 261 398
rect 261 397 262 398
rect 262 397 263 398
rect 263 397 264 398
rect 264 397 265 398
rect 265 397 266 398
rect 266 397 267 398
rect 267 397 268 398
rect 268 397 269 398
rect 269 397 270 398
rect 270 397 271 398
rect 271 397 272 398
rect 272 397 273 398
rect 273 397 274 398
rect 274 397 275 398
rect 481 397 482 398
rect 482 397 483 398
rect 483 397 484 398
rect 484 397 485 398
rect 485 397 486 398
rect 486 397 487 398
rect 487 397 488 398
rect 488 397 489 398
rect 489 397 490 398
rect 75 396 76 397
rect 76 396 77 397
rect 77 396 78 397
rect 78 396 79 397
rect 79 396 80 397
rect 80 396 81 397
rect 81 396 82 397
rect 82 396 83 397
rect 83 396 84 397
rect 84 396 85 397
rect 85 396 86 397
rect 119 396 120 397
rect 120 396 121 397
rect 121 396 122 397
rect 122 396 123 397
rect 123 396 124 397
rect 124 396 125 397
rect 125 396 126 397
rect 126 396 127 397
rect 203 396 204 397
rect 204 396 205 397
rect 205 396 206 397
rect 206 396 207 397
rect 207 396 208 397
rect 208 396 209 397
rect 209 396 210 397
rect 210 396 211 397
rect 211 396 212 397
rect 212 396 213 397
rect 226 396 227 397
rect 227 396 228 397
rect 228 396 229 397
rect 229 396 230 397
rect 230 396 231 397
rect 231 396 232 397
rect 232 396 233 397
rect 233 396 234 397
rect 234 396 235 397
rect 235 396 236 397
rect 236 396 237 397
rect 237 396 238 397
rect 238 396 239 397
rect 239 396 240 397
rect 240 396 241 397
rect 241 396 242 397
rect 242 396 243 397
rect 243 396 244 397
rect 244 396 245 397
rect 245 396 246 397
rect 246 396 247 397
rect 247 396 248 397
rect 248 396 249 397
rect 249 396 250 397
rect 250 396 251 397
rect 251 396 252 397
rect 252 396 253 397
rect 253 396 254 397
rect 254 396 255 397
rect 255 396 256 397
rect 256 396 257 397
rect 257 396 258 397
rect 258 396 259 397
rect 259 396 260 397
rect 260 396 261 397
rect 261 396 262 397
rect 262 396 263 397
rect 263 396 264 397
rect 264 396 265 397
rect 265 396 266 397
rect 266 396 267 397
rect 267 396 268 397
rect 268 396 269 397
rect 269 396 270 397
rect 270 396 271 397
rect 271 396 272 397
rect 272 396 273 397
rect 273 396 274 397
rect 274 396 275 397
rect 275 396 276 397
rect 276 396 277 397
rect 481 396 482 397
rect 482 396 483 397
rect 483 396 484 397
rect 484 396 485 397
rect 485 396 486 397
rect 486 396 487 397
rect 487 396 488 397
rect 488 396 489 397
rect 489 396 490 397
rect 74 395 75 396
rect 75 395 76 396
rect 76 395 77 396
rect 77 395 78 396
rect 78 395 79 396
rect 79 395 80 396
rect 80 395 81 396
rect 81 395 82 396
rect 82 395 83 396
rect 83 395 84 396
rect 84 395 85 396
rect 118 395 119 396
rect 119 395 120 396
rect 120 395 121 396
rect 121 395 122 396
rect 122 395 123 396
rect 123 395 124 396
rect 202 395 203 396
rect 203 395 204 396
rect 204 395 205 396
rect 205 395 206 396
rect 206 395 207 396
rect 207 395 208 396
rect 208 395 209 396
rect 209 395 210 396
rect 223 395 224 396
rect 224 395 225 396
rect 225 395 226 396
rect 226 395 227 396
rect 227 395 228 396
rect 228 395 229 396
rect 229 395 230 396
rect 230 395 231 396
rect 231 395 232 396
rect 232 395 233 396
rect 233 395 234 396
rect 234 395 235 396
rect 235 395 236 396
rect 236 395 237 396
rect 237 395 238 396
rect 238 395 239 396
rect 239 395 240 396
rect 240 395 241 396
rect 241 395 242 396
rect 242 395 243 396
rect 243 395 244 396
rect 244 395 245 396
rect 245 395 246 396
rect 246 395 247 396
rect 247 395 248 396
rect 248 395 249 396
rect 249 395 250 396
rect 250 395 251 396
rect 251 395 252 396
rect 252 395 253 396
rect 253 395 254 396
rect 254 395 255 396
rect 255 395 256 396
rect 256 395 257 396
rect 257 395 258 396
rect 258 395 259 396
rect 259 395 260 396
rect 260 395 261 396
rect 261 395 262 396
rect 262 395 263 396
rect 263 395 264 396
rect 264 395 265 396
rect 265 395 266 396
rect 266 395 267 396
rect 267 395 268 396
rect 268 395 269 396
rect 269 395 270 396
rect 270 395 271 396
rect 271 395 272 396
rect 272 395 273 396
rect 273 395 274 396
rect 274 395 275 396
rect 275 395 276 396
rect 276 395 277 396
rect 277 395 278 396
rect 278 395 279 396
rect 482 395 483 396
rect 483 395 484 396
rect 484 395 485 396
rect 485 395 486 396
rect 486 395 487 396
rect 487 395 488 396
rect 488 395 489 396
rect 489 395 490 396
rect 490 395 491 396
rect 73 394 74 395
rect 74 394 75 395
rect 75 394 76 395
rect 76 394 77 395
rect 77 394 78 395
rect 78 394 79 395
rect 79 394 80 395
rect 80 394 81 395
rect 81 394 82 395
rect 82 394 83 395
rect 83 394 84 395
rect 201 394 202 395
rect 202 394 203 395
rect 203 394 204 395
rect 204 394 205 395
rect 205 394 206 395
rect 206 394 207 395
rect 207 394 208 395
rect 221 394 222 395
rect 222 394 223 395
rect 223 394 224 395
rect 224 394 225 395
rect 225 394 226 395
rect 226 394 227 395
rect 227 394 228 395
rect 228 394 229 395
rect 229 394 230 395
rect 230 394 231 395
rect 231 394 232 395
rect 232 394 233 395
rect 233 394 234 395
rect 234 394 235 395
rect 235 394 236 395
rect 236 394 237 395
rect 237 394 238 395
rect 238 394 239 395
rect 239 394 240 395
rect 240 394 241 395
rect 241 394 242 395
rect 242 394 243 395
rect 243 394 244 395
rect 244 394 245 395
rect 245 394 246 395
rect 246 394 247 395
rect 247 394 248 395
rect 248 394 249 395
rect 249 394 250 395
rect 250 394 251 395
rect 251 394 252 395
rect 252 394 253 395
rect 253 394 254 395
rect 254 394 255 395
rect 255 394 256 395
rect 256 394 257 395
rect 257 394 258 395
rect 258 394 259 395
rect 259 394 260 395
rect 260 394 261 395
rect 261 394 262 395
rect 262 394 263 395
rect 263 394 264 395
rect 264 394 265 395
rect 265 394 266 395
rect 266 394 267 395
rect 267 394 268 395
rect 268 394 269 395
rect 269 394 270 395
rect 270 394 271 395
rect 271 394 272 395
rect 272 394 273 395
rect 273 394 274 395
rect 274 394 275 395
rect 275 394 276 395
rect 276 394 277 395
rect 277 394 278 395
rect 278 394 279 395
rect 279 394 280 395
rect 280 394 281 395
rect 482 394 483 395
rect 483 394 484 395
rect 484 394 485 395
rect 485 394 486 395
rect 486 394 487 395
rect 487 394 488 395
rect 488 394 489 395
rect 489 394 490 395
rect 490 394 491 395
rect 73 393 74 394
rect 74 393 75 394
rect 75 393 76 394
rect 76 393 77 394
rect 77 393 78 394
rect 78 393 79 394
rect 79 393 80 394
rect 80 393 81 394
rect 81 393 82 394
rect 82 393 83 394
rect 83 393 84 394
rect 201 393 202 394
rect 202 393 203 394
rect 203 393 204 394
rect 204 393 205 394
rect 205 393 206 394
rect 218 393 219 394
rect 219 393 220 394
rect 220 393 221 394
rect 221 393 222 394
rect 222 393 223 394
rect 223 393 224 394
rect 224 393 225 394
rect 225 393 226 394
rect 226 393 227 394
rect 227 393 228 394
rect 228 393 229 394
rect 229 393 230 394
rect 230 393 231 394
rect 231 393 232 394
rect 232 393 233 394
rect 233 393 234 394
rect 234 393 235 394
rect 235 393 236 394
rect 236 393 237 394
rect 237 393 238 394
rect 238 393 239 394
rect 239 393 240 394
rect 240 393 241 394
rect 241 393 242 394
rect 242 393 243 394
rect 243 393 244 394
rect 244 393 245 394
rect 245 393 246 394
rect 246 393 247 394
rect 247 393 248 394
rect 248 393 249 394
rect 249 393 250 394
rect 250 393 251 394
rect 251 393 252 394
rect 252 393 253 394
rect 253 393 254 394
rect 254 393 255 394
rect 255 393 256 394
rect 256 393 257 394
rect 257 393 258 394
rect 258 393 259 394
rect 259 393 260 394
rect 260 393 261 394
rect 261 393 262 394
rect 262 393 263 394
rect 263 393 264 394
rect 264 393 265 394
rect 265 393 266 394
rect 266 393 267 394
rect 267 393 268 394
rect 268 393 269 394
rect 269 393 270 394
rect 270 393 271 394
rect 271 393 272 394
rect 272 393 273 394
rect 273 393 274 394
rect 274 393 275 394
rect 275 393 276 394
rect 276 393 277 394
rect 277 393 278 394
rect 278 393 279 394
rect 279 393 280 394
rect 280 393 281 394
rect 281 393 282 394
rect 282 393 283 394
rect 283 393 284 394
rect 482 393 483 394
rect 483 393 484 394
rect 484 393 485 394
rect 485 393 486 394
rect 486 393 487 394
rect 487 393 488 394
rect 488 393 489 394
rect 489 393 490 394
rect 490 393 491 394
rect 72 392 73 393
rect 73 392 74 393
rect 74 392 75 393
rect 75 392 76 393
rect 76 392 77 393
rect 77 392 78 393
rect 78 392 79 393
rect 79 392 80 393
rect 80 392 81 393
rect 81 392 82 393
rect 82 392 83 393
rect 200 392 201 393
rect 201 392 202 393
rect 202 392 203 393
rect 203 392 204 393
rect 216 392 217 393
rect 217 392 218 393
rect 218 392 219 393
rect 219 392 220 393
rect 220 392 221 393
rect 221 392 222 393
rect 222 392 223 393
rect 223 392 224 393
rect 224 392 225 393
rect 225 392 226 393
rect 226 392 227 393
rect 227 392 228 393
rect 228 392 229 393
rect 229 392 230 393
rect 230 392 231 393
rect 231 392 232 393
rect 232 392 233 393
rect 233 392 234 393
rect 234 392 235 393
rect 235 392 236 393
rect 236 392 237 393
rect 237 392 238 393
rect 238 392 239 393
rect 239 392 240 393
rect 240 392 241 393
rect 241 392 242 393
rect 242 392 243 393
rect 243 392 244 393
rect 244 392 245 393
rect 245 392 246 393
rect 246 392 247 393
rect 247 392 248 393
rect 248 392 249 393
rect 249 392 250 393
rect 250 392 251 393
rect 251 392 252 393
rect 252 392 253 393
rect 253 392 254 393
rect 254 392 255 393
rect 255 392 256 393
rect 256 392 257 393
rect 257 392 258 393
rect 258 392 259 393
rect 259 392 260 393
rect 260 392 261 393
rect 261 392 262 393
rect 262 392 263 393
rect 263 392 264 393
rect 264 392 265 393
rect 265 392 266 393
rect 266 392 267 393
rect 267 392 268 393
rect 268 392 269 393
rect 269 392 270 393
rect 270 392 271 393
rect 271 392 272 393
rect 272 392 273 393
rect 273 392 274 393
rect 274 392 275 393
rect 275 392 276 393
rect 276 392 277 393
rect 277 392 278 393
rect 278 392 279 393
rect 279 392 280 393
rect 280 392 281 393
rect 281 392 282 393
rect 282 392 283 393
rect 283 392 284 393
rect 284 392 285 393
rect 285 392 286 393
rect 286 392 287 393
rect 287 392 288 393
rect 288 392 289 393
rect 289 392 290 393
rect 483 392 484 393
rect 484 392 485 393
rect 485 392 486 393
rect 486 392 487 393
rect 487 392 488 393
rect 488 392 489 393
rect 489 392 490 393
rect 490 392 491 393
rect 491 392 492 393
rect 71 391 72 392
rect 72 391 73 392
rect 73 391 74 392
rect 74 391 75 392
rect 75 391 76 392
rect 76 391 77 392
rect 77 391 78 392
rect 78 391 79 392
rect 79 391 80 392
rect 80 391 81 392
rect 81 391 82 392
rect 199 391 200 392
rect 200 391 201 392
rect 201 391 202 392
rect 214 391 215 392
rect 215 391 216 392
rect 216 391 217 392
rect 217 391 218 392
rect 218 391 219 392
rect 219 391 220 392
rect 220 391 221 392
rect 221 391 222 392
rect 222 391 223 392
rect 223 391 224 392
rect 224 391 225 392
rect 225 391 226 392
rect 226 391 227 392
rect 227 391 228 392
rect 228 391 229 392
rect 229 391 230 392
rect 230 391 231 392
rect 231 391 232 392
rect 232 391 233 392
rect 233 391 234 392
rect 234 391 235 392
rect 235 391 236 392
rect 236 391 237 392
rect 237 391 238 392
rect 238 391 239 392
rect 239 391 240 392
rect 240 391 241 392
rect 241 391 242 392
rect 242 391 243 392
rect 243 391 244 392
rect 244 391 245 392
rect 245 391 246 392
rect 246 391 247 392
rect 247 391 248 392
rect 248 391 249 392
rect 249 391 250 392
rect 250 391 251 392
rect 251 391 252 392
rect 252 391 253 392
rect 253 391 254 392
rect 254 391 255 392
rect 255 391 256 392
rect 256 391 257 392
rect 257 391 258 392
rect 258 391 259 392
rect 259 391 260 392
rect 260 391 261 392
rect 261 391 262 392
rect 262 391 263 392
rect 263 391 264 392
rect 264 391 265 392
rect 265 391 266 392
rect 266 391 267 392
rect 267 391 268 392
rect 268 391 269 392
rect 269 391 270 392
rect 270 391 271 392
rect 271 391 272 392
rect 272 391 273 392
rect 273 391 274 392
rect 274 391 275 392
rect 275 391 276 392
rect 276 391 277 392
rect 277 391 278 392
rect 278 391 279 392
rect 279 391 280 392
rect 280 391 281 392
rect 281 391 282 392
rect 282 391 283 392
rect 283 391 284 392
rect 284 391 285 392
rect 285 391 286 392
rect 286 391 287 392
rect 287 391 288 392
rect 288 391 289 392
rect 289 391 290 392
rect 290 391 291 392
rect 291 391 292 392
rect 292 391 293 392
rect 293 391 294 392
rect 294 391 295 392
rect 295 391 296 392
rect 483 391 484 392
rect 484 391 485 392
rect 485 391 486 392
rect 486 391 487 392
rect 487 391 488 392
rect 488 391 489 392
rect 489 391 490 392
rect 490 391 491 392
rect 491 391 492 392
rect 71 390 72 391
rect 72 390 73 391
rect 73 390 74 391
rect 74 390 75 391
rect 75 390 76 391
rect 76 390 77 391
rect 77 390 78 391
rect 78 390 79 391
rect 79 390 80 391
rect 80 390 81 391
rect 199 390 200 391
rect 212 390 213 391
rect 213 390 214 391
rect 214 390 215 391
rect 215 390 216 391
rect 216 390 217 391
rect 217 390 218 391
rect 218 390 219 391
rect 219 390 220 391
rect 220 390 221 391
rect 221 390 222 391
rect 222 390 223 391
rect 223 390 224 391
rect 224 390 225 391
rect 225 390 226 391
rect 226 390 227 391
rect 227 390 228 391
rect 228 390 229 391
rect 229 390 230 391
rect 230 390 231 391
rect 231 390 232 391
rect 232 390 233 391
rect 233 390 234 391
rect 234 390 235 391
rect 235 390 236 391
rect 236 390 237 391
rect 237 390 238 391
rect 238 390 239 391
rect 239 390 240 391
rect 240 390 241 391
rect 241 390 242 391
rect 242 390 243 391
rect 243 390 244 391
rect 244 390 245 391
rect 245 390 246 391
rect 246 390 247 391
rect 247 390 248 391
rect 248 390 249 391
rect 249 390 250 391
rect 250 390 251 391
rect 251 390 252 391
rect 252 390 253 391
rect 253 390 254 391
rect 254 390 255 391
rect 255 390 256 391
rect 256 390 257 391
rect 257 390 258 391
rect 258 390 259 391
rect 259 390 260 391
rect 260 390 261 391
rect 261 390 262 391
rect 262 390 263 391
rect 263 390 264 391
rect 264 390 265 391
rect 265 390 266 391
rect 266 390 267 391
rect 267 390 268 391
rect 268 390 269 391
rect 269 390 270 391
rect 270 390 271 391
rect 271 390 272 391
rect 272 390 273 391
rect 273 390 274 391
rect 274 390 275 391
rect 275 390 276 391
rect 276 390 277 391
rect 277 390 278 391
rect 278 390 279 391
rect 279 390 280 391
rect 280 390 281 391
rect 281 390 282 391
rect 282 390 283 391
rect 283 390 284 391
rect 284 390 285 391
rect 285 390 286 391
rect 286 390 287 391
rect 287 390 288 391
rect 288 390 289 391
rect 289 390 290 391
rect 290 390 291 391
rect 291 390 292 391
rect 292 390 293 391
rect 293 390 294 391
rect 294 390 295 391
rect 295 390 296 391
rect 296 390 297 391
rect 297 390 298 391
rect 298 390 299 391
rect 299 390 300 391
rect 300 390 301 391
rect 483 390 484 391
rect 484 390 485 391
rect 485 390 486 391
rect 486 390 487 391
rect 487 390 488 391
rect 488 390 489 391
rect 489 390 490 391
rect 490 390 491 391
rect 491 390 492 391
rect 70 389 71 390
rect 71 389 72 390
rect 72 389 73 390
rect 73 389 74 390
rect 74 389 75 390
rect 75 389 76 390
rect 76 389 77 390
rect 77 389 78 390
rect 78 389 79 390
rect 79 389 80 390
rect 80 389 81 390
rect 211 389 212 390
rect 212 389 213 390
rect 213 389 214 390
rect 214 389 215 390
rect 215 389 216 390
rect 216 389 217 390
rect 217 389 218 390
rect 218 389 219 390
rect 219 389 220 390
rect 220 389 221 390
rect 221 389 222 390
rect 222 389 223 390
rect 223 389 224 390
rect 224 389 225 390
rect 225 389 226 390
rect 226 389 227 390
rect 227 389 228 390
rect 228 389 229 390
rect 229 389 230 390
rect 230 389 231 390
rect 231 389 232 390
rect 232 389 233 390
rect 233 389 234 390
rect 234 389 235 390
rect 235 389 236 390
rect 236 389 237 390
rect 237 389 238 390
rect 238 389 239 390
rect 239 389 240 390
rect 240 389 241 390
rect 241 389 242 390
rect 242 389 243 390
rect 243 389 244 390
rect 244 389 245 390
rect 245 389 246 390
rect 246 389 247 390
rect 247 389 248 390
rect 248 389 249 390
rect 249 389 250 390
rect 250 389 251 390
rect 251 389 252 390
rect 252 389 253 390
rect 253 389 254 390
rect 254 389 255 390
rect 255 389 256 390
rect 256 389 257 390
rect 257 389 258 390
rect 258 389 259 390
rect 259 389 260 390
rect 260 389 261 390
rect 261 389 262 390
rect 262 389 263 390
rect 263 389 264 390
rect 264 389 265 390
rect 265 389 266 390
rect 266 389 267 390
rect 267 389 268 390
rect 268 389 269 390
rect 269 389 270 390
rect 270 389 271 390
rect 271 389 272 390
rect 272 389 273 390
rect 273 389 274 390
rect 274 389 275 390
rect 275 389 276 390
rect 276 389 277 390
rect 277 389 278 390
rect 278 389 279 390
rect 279 389 280 390
rect 280 389 281 390
rect 281 389 282 390
rect 282 389 283 390
rect 283 389 284 390
rect 284 389 285 390
rect 285 389 286 390
rect 286 389 287 390
rect 287 389 288 390
rect 288 389 289 390
rect 289 389 290 390
rect 290 389 291 390
rect 291 389 292 390
rect 292 389 293 390
rect 293 389 294 390
rect 294 389 295 390
rect 295 389 296 390
rect 296 389 297 390
rect 297 389 298 390
rect 298 389 299 390
rect 299 389 300 390
rect 300 389 301 390
rect 301 389 302 390
rect 302 389 303 390
rect 303 389 304 390
rect 304 389 305 390
rect 483 389 484 390
rect 484 389 485 390
rect 485 389 486 390
rect 486 389 487 390
rect 487 389 488 390
rect 488 389 489 390
rect 489 389 490 390
rect 490 389 491 390
rect 491 389 492 390
rect 69 388 70 389
rect 70 388 71 389
rect 71 388 72 389
rect 72 388 73 389
rect 73 388 74 389
rect 74 388 75 389
rect 75 388 76 389
rect 76 388 77 389
rect 77 388 78 389
rect 78 388 79 389
rect 79 388 80 389
rect 209 388 210 389
rect 210 388 211 389
rect 211 388 212 389
rect 212 388 213 389
rect 213 388 214 389
rect 214 388 215 389
rect 215 388 216 389
rect 216 388 217 389
rect 217 388 218 389
rect 218 388 219 389
rect 219 388 220 389
rect 220 388 221 389
rect 221 388 222 389
rect 222 388 223 389
rect 223 388 224 389
rect 224 388 225 389
rect 225 388 226 389
rect 226 388 227 389
rect 227 388 228 389
rect 228 388 229 389
rect 229 388 230 389
rect 230 388 231 389
rect 231 388 232 389
rect 232 388 233 389
rect 233 388 234 389
rect 234 388 235 389
rect 235 388 236 389
rect 236 388 237 389
rect 237 388 238 389
rect 238 388 239 389
rect 239 388 240 389
rect 240 388 241 389
rect 241 388 242 389
rect 242 388 243 389
rect 243 388 244 389
rect 244 388 245 389
rect 245 388 246 389
rect 246 388 247 389
rect 247 388 248 389
rect 248 388 249 389
rect 249 388 250 389
rect 250 388 251 389
rect 251 388 252 389
rect 252 388 253 389
rect 253 388 254 389
rect 254 388 255 389
rect 255 388 256 389
rect 256 388 257 389
rect 257 388 258 389
rect 258 388 259 389
rect 259 388 260 389
rect 260 388 261 389
rect 261 388 262 389
rect 262 388 263 389
rect 263 388 264 389
rect 264 388 265 389
rect 265 388 266 389
rect 266 388 267 389
rect 267 388 268 389
rect 268 388 269 389
rect 269 388 270 389
rect 270 388 271 389
rect 271 388 272 389
rect 272 388 273 389
rect 273 388 274 389
rect 274 388 275 389
rect 275 388 276 389
rect 276 388 277 389
rect 277 388 278 389
rect 278 388 279 389
rect 279 388 280 389
rect 280 388 281 389
rect 281 388 282 389
rect 282 388 283 389
rect 283 388 284 389
rect 284 388 285 389
rect 285 388 286 389
rect 286 388 287 389
rect 287 388 288 389
rect 288 388 289 389
rect 289 388 290 389
rect 290 388 291 389
rect 291 388 292 389
rect 292 388 293 389
rect 293 388 294 389
rect 294 388 295 389
rect 295 388 296 389
rect 296 388 297 389
rect 297 388 298 389
rect 298 388 299 389
rect 299 388 300 389
rect 300 388 301 389
rect 301 388 302 389
rect 302 388 303 389
rect 303 388 304 389
rect 304 388 305 389
rect 305 388 306 389
rect 306 388 307 389
rect 484 388 485 389
rect 485 388 486 389
rect 486 388 487 389
rect 487 388 488 389
rect 488 388 489 389
rect 489 388 490 389
rect 490 388 491 389
rect 491 388 492 389
rect 69 387 70 388
rect 70 387 71 388
rect 71 387 72 388
rect 72 387 73 388
rect 73 387 74 388
rect 74 387 75 388
rect 75 387 76 388
rect 76 387 77 388
rect 77 387 78 388
rect 78 387 79 388
rect 208 387 209 388
rect 209 387 210 388
rect 210 387 211 388
rect 211 387 212 388
rect 212 387 213 388
rect 213 387 214 388
rect 214 387 215 388
rect 215 387 216 388
rect 216 387 217 388
rect 217 387 218 388
rect 218 387 219 388
rect 219 387 220 388
rect 220 387 221 388
rect 221 387 222 388
rect 222 387 223 388
rect 223 387 224 388
rect 224 387 225 388
rect 225 387 226 388
rect 226 387 227 388
rect 227 387 228 388
rect 228 387 229 388
rect 229 387 230 388
rect 230 387 231 388
rect 231 387 232 388
rect 232 387 233 388
rect 233 387 234 388
rect 234 387 235 388
rect 235 387 236 388
rect 236 387 237 388
rect 237 387 238 388
rect 238 387 239 388
rect 239 387 240 388
rect 240 387 241 388
rect 241 387 242 388
rect 242 387 243 388
rect 243 387 244 388
rect 244 387 245 388
rect 245 387 246 388
rect 246 387 247 388
rect 247 387 248 388
rect 248 387 249 388
rect 249 387 250 388
rect 250 387 251 388
rect 251 387 252 388
rect 252 387 253 388
rect 253 387 254 388
rect 254 387 255 388
rect 255 387 256 388
rect 256 387 257 388
rect 257 387 258 388
rect 258 387 259 388
rect 259 387 260 388
rect 260 387 261 388
rect 261 387 262 388
rect 262 387 263 388
rect 263 387 264 388
rect 264 387 265 388
rect 265 387 266 388
rect 266 387 267 388
rect 267 387 268 388
rect 268 387 269 388
rect 269 387 270 388
rect 270 387 271 388
rect 271 387 272 388
rect 272 387 273 388
rect 273 387 274 388
rect 274 387 275 388
rect 275 387 276 388
rect 276 387 277 388
rect 277 387 278 388
rect 278 387 279 388
rect 279 387 280 388
rect 280 387 281 388
rect 281 387 282 388
rect 282 387 283 388
rect 283 387 284 388
rect 284 387 285 388
rect 285 387 286 388
rect 286 387 287 388
rect 287 387 288 388
rect 288 387 289 388
rect 289 387 290 388
rect 290 387 291 388
rect 291 387 292 388
rect 292 387 293 388
rect 293 387 294 388
rect 294 387 295 388
rect 295 387 296 388
rect 296 387 297 388
rect 297 387 298 388
rect 298 387 299 388
rect 299 387 300 388
rect 300 387 301 388
rect 301 387 302 388
rect 302 387 303 388
rect 303 387 304 388
rect 304 387 305 388
rect 305 387 306 388
rect 306 387 307 388
rect 307 387 308 388
rect 308 387 309 388
rect 309 387 310 388
rect 484 387 485 388
rect 485 387 486 388
rect 486 387 487 388
rect 487 387 488 388
rect 488 387 489 388
rect 489 387 490 388
rect 490 387 491 388
rect 491 387 492 388
rect 492 387 493 388
rect 68 386 69 387
rect 69 386 70 387
rect 70 386 71 387
rect 71 386 72 387
rect 72 386 73 387
rect 73 386 74 387
rect 74 386 75 387
rect 75 386 76 387
rect 76 386 77 387
rect 77 386 78 387
rect 78 386 79 387
rect 207 386 208 387
rect 208 386 209 387
rect 209 386 210 387
rect 210 386 211 387
rect 211 386 212 387
rect 212 386 213 387
rect 213 386 214 387
rect 214 386 215 387
rect 215 386 216 387
rect 216 386 217 387
rect 217 386 218 387
rect 218 386 219 387
rect 219 386 220 387
rect 220 386 221 387
rect 221 386 222 387
rect 222 386 223 387
rect 223 386 224 387
rect 224 386 225 387
rect 225 386 226 387
rect 226 386 227 387
rect 227 386 228 387
rect 228 386 229 387
rect 229 386 230 387
rect 230 386 231 387
rect 231 386 232 387
rect 232 386 233 387
rect 233 386 234 387
rect 234 386 235 387
rect 235 386 236 387
rect 236 386 237 387
rect 237 386 238 387
rect 238 386 239 387
rect 239 386 240 387
rect 240 386 241 387
rect 241 386 242 387
rect 242 386 243 387
rect 243 386 244 387
rect 244 386 245 387
rect 245 386 246 387
rect 246 386 247 387
rect 247 386 248 387
rect 248 386 249 387
rect 249 386 250 387
rect 250 386 251 387
rect 251 386 252 387
rect 252 386 253 387
rect 253 386 254 387
rect 254 386 255 387
rect 255 386 256 387
rect 256 386 257 387
rect 257 386 258 387
rect 258 386 259 387
rect 259 386 260 387
rect 260 386 261 387
rect 261 386 262 387
rect 262 386 263 387
rect 263 386 264 387
rect 264 386 265 387
rect 265 386 266 387
rect 266 386 267 387
rect 267 386 268 387
rect 268 386 269 387
rect 269 386 270 387
rect 270 386 271 387
rect 271 386 272 387
rect 272 386 273 387
rect 273 386 274 387
rect 274 386 275 387
rect 275 386 276 387
rect 276 386 277 387
rect 277 386 278 387
rect 278 386 279 387
rect 279 386 280 387
rect 280 386 281 387
rect 281 386 282 387
rect 282 386 283 387
rect 283 386 284 387
rect 284 386 285 387
rect 285 386 286 387
rect 286 386 287 387
rect 287 386 288 387
rect 288 386 289 387
rect 289 386 290 387
rect 290 386 291 387
rect 291 386 292 387
rect 292 386 293 387
rect 293 386 294 387
rect 294 386 295 387
rect 295 386 296 387
rect 296 386 297 387
rect 297 386 298 387
rect 298 386 299 387
rect 299 386 300 387
rect 300 386 301 387
rect 301 386 302 387
rect 302 386 303 387
rect 303 386 304 387
rect 304 386 305 387
rect 305 386 306 387
rect 306 386 307 387
rect 307 386 308 387
rect 308 386 309 387
rect 309 386 310 387
rect 310 386 311 387
rect 311 386 312 387
rect 484 386 485 387
rect 485 386 486 387
rect 486 386 487 387
rect 487 386 488 387
rect 488 386 489 387
rect 489 386 490 387
rect 490 386 491 387
rect 491 386 492 387
rect 492 386 493 387
rect 68 385 69 386
rect 69 385 70 386
rect 70 385 71 386
rect 71 385 72 386
rect 72 385 73 386
rect 73 385 74 386
rect 74 385 75 386
rect 75 385 76 386
rect 76 385 77 386
rect 77 385 78 386
rect 205 385 206 386
rect 206 385 207 386
rect 207 385 208 386
rect 208 385 209 386
rect 209 385 210 386
rect 210 385 211 386
rect 211 385 212 386
rect 212 385 213 386
rect 213 385 214 386
rect 214 385 215 386
rect 215 385 216 386
rect 216 385 217 386
rect 217 385 218 386
rect 218 385 219 386
rect 219 385 220 386
rect 220 385 221 386
rect 221 385 222 386
rect 222 385 223 386
rect 223 385 224 386
rect 224 385 225 386
rect 225 385 226 386
rect 226 385 227 386
rect 227 385 228 386
rect 228 385 229 386
rect 229 385 230 386
rect 230 385 231 386
rect 231 385 232 386
rect 232 385 233 386
rect 233 385 234 386
rect 234 385 235 386
rect 235 385 236 386
rect 236 385 237 386
rect 237 385 238 386
rect 238 385 239 386
rect 239 385 240 386
rect 240 385 241 386
rect 241 385 242 386
rect 242 385 243 386
rect 243 385 244 386
rect 244 385 245 386
rect 245 385 246 386
rect 246 385 247 386
rect 247 385 248 386
rect 248 385 249 386
rect 249 385 250 386
rect 250 385 251 386
rect 251 385 252 386
rect 252 385 253 386
rect 253 385 254 386
rect 254 385 255 386
rect 255 385 256 386
rect 256 385 257 386
rect 257 385 258 386
rect 258 385 259 386
rect 259 385 260 386
rect 260 385 261 386
rect 261 385 262 386
rect 262 385 263 386
rect 263 385 264 386
rect 264 385 265 386
rect 265 385 266 386
rect 266 385 267 386
rect 267 385 268 386
rect 268 385 269 386
rect 269 385 270 386
rect 270 385 271 386
rect 271 385 272 386
rect 272 385 273 386
rect 273 385 274 386
rect 274 385 275 386
rect 275 385 276 386
rect 276 385 277 386
rect 277 385 278 386
rect 278 385 279 386
rect 279 385 280 386
rect 280 385 281 386
rect 281 385 282 386
rect 282 385 283 386
rect 283 385 284 386
rect 284 385 285 386
rect 285 385 286 386
rect 286 385 287 386
rect 287 385 288 386
rect 288 385 289 386
rect 289 385 290 386
rect 290 385 291 386
rect 291 385 292 386
rect 292 385 293 386
rect 293 385 294 386
rect 294 385 295 386
rect 295 385 296 386
rect 296 385 297 386
rect 297 385 298 386
rect 298 385 299 386
rect 299 385 300 386
rect 300 385 301 386
rect 301 385 302 386
rect 302 385 303 386
rect 303 385 304 386
rect 304 385 305 386
rect 305 385 306 386
rect 306 385 307 386
rect 307 385 308 386
rect 308 385 309 386
rect 309 385 310 386
rect 310 385 311 386
rect 311 385 312 386
rect 312 385 313 386
rect 313 385 314 386
rect 314 385 315 386
rect 484 385 485 386
rect 485 385 486 386
rect 486 385 487 386
rect 487 385 488 386
rect 488 385 489 386
rect 489 385 490 386
rect 490 385 491 386
rect 491 385 492 386
rect 492 385 493 386
rect 67 384 68 385
rect 68 384 69 385
rect 69 384 70 385
rect 70 384 71 385
rect 71 384 72 385
rect 72 384 73 385
rect 73 384 74 385
rect 74 384 75 385
rect 75 384 76 385
rect 76 384 77 385
rect 204 384 205 385
rect 205 384 206 385
rect 206 384 207 385
rect 207 384 208 385
rect 208 384 209 385
rect 209 384 210 385
rect 210 384 211 385
rect 211 384 212 385
rect 212 384 213 385
rect 213 384 214 385
rect 214 384 215 385
rect 215 384 216 385
rect 216 384 217 385
rect 217 384 218 385
rect 218 384 219 385
rect 219 384 220 385
rect 220 384 221 385
rect 221 384 222 385
rect 222 384 223 385
rect 223 384 224 385
rect 224 384 225 385
rect 225 384 226 385
rect 226 384 227 385
rect 227 384 228 385
rect 228 384 229 385
rect 229 384 230 385
rect 230 384 231 385
rect 231 384 232 385
rect 232 384 233 385
rect 233 384 234 385
rect 234 384 235 385
rect 235 384 236 385
rect 236 384 237 385
rect 237 384 238 385
rect 238 384 239 385
rect 239 384 240 385
rect 240 384 241 385
rect 241 384 242 385
rect 242 384 243 385
rect 243 384 244 385
rect 244 384 245 385
rect 245 384 246 385
rect 246 384 247 385
rect 247 384 248 385
rect 248 384 249 385
rect 249 384 250 385
rect 250 384 251 385
rect 251 384 252 385
rect 252 384 253 385
rect 253 384 254 385
rect 254 384 255 385
rect 255 384 256 385
rect 256 384 257 385
rect 257 384 258 385
rect 258 384 259 385
rect 259 384 260 385
rect 260 384 261 385
rect 261 384 262 385
rect 262 384 263 385
rect 263 384 264 385
rect 264 384 265 385
rect 265 384 266 385
rect 266 384 267 385
rect 267 384 268 385
rect 268 384 269 385
rect 269 384 270 385
rect 270 384 271 385
rect 271 384 272 385
rect 272 384 273 385
rect 273 384 274 385
rect 274 384 275 385
rect 275 384 276 385
rect 276 384 277 385
rect 277 384 278 385
rect 278 384 279 385
rect 279 384 280 385
rect 280 384 281 385
rect 281 384 282 385
rect 282 384 283 385
rect 283 384 284 385
rect 284 384 285 385
rect 285 384 286 385
rect 286 384 287 385
rect 287 384 288 385
rect 288 384 289 385
rect 289 384 290 385
rect 290 384 291 385
rect 291 384 292 385
rect 292 384 293 385
rect 293 384 294 385
rect 294 384 295 385
rect 295 384 296 385
rect 296 384 297 385
rect 297 384 298 385
rect 298 384 299 385
rect 299 384 300 385
rect 300 384 301 385
rect 301 384 302 385
rect 302 384 303 385
rect 303 384 304 385
rect 304 384 305 385
rect 305 384 306 385
rect 306 384 307 385
rect 307 384 308 385
rect 308 384 309 385
rect 309 384 310 385
rect 310 384 311 385
rect 311 384 312 385
rect 312 384 313 385
rect 313 384 314 385
rect 314 384 315 385
rect 315 384 316 385
rect 484 384 485 385
rect 485 384 486 385
rect 486 384 487 385
rect 487 384 488 385
rect 488 384 489 385
rect 489 384 490 385
rect 490 384 491 385
rect 491 384 492 385
rect 492 384 493 385
rect 67 383 68 384
rect 68 383 69 384
rect 69 383 70 384
rect 70 383 71 384
rect 71 383 72 384
rect 72 383 73 384
rect 73 383 74 384
rect 74 383 75 384
rect 75 383 76 384
rect 76 383 77 384
rect 203 383 204 384
rect 204 383 205 384
rect 205 383 206 384
rect 206 383 207 384
rect 207 383 208 384
rect 208 383 209 384
rect 209 383 210 384
rect 210 383 211 384
rect 211 383 212 384
rect 212 383 213 384
rect 213 383 214 384
rect 214 383 215 384
rect 215 383 216 384
rect 216 383 217 384
rect 217 383 218 384
rect 218 383 219 384
rect 219 383 220 384
rect 220 383 221 384
rect 221 383 222 384
rect 222 383 223 384
rect 223 383 224 384
rect 224 383 225 384
rect 225 383 226 384
rect 226 383 227 384
rect 227 383 228 384
rect 228 383 229 384
rect 229 383 230 384
rect 230 383 231 384
rect 231 383 232 384
rect 232 383 233 384
rect 233 383 234 384
rect 234 383 235 384
rect 235 383 236 384
rect 236 383 237 384
rect 237 383 238 384
rect 238 383 239 384
rect 239 383 240 384
rect 240 383 241 384
rect 241 383 242 384
rect 242 383 243 384
rect 243 383 244 384
rect 244 383 245 384
rect 245 383 246 384
rect 246 383 247 384
rect 247 383 248 384
rect 248 383 249 384
rect 249 383 250 384
rect 250 383 251 384
rect 251 383 252 384
rect 252 383 253 384
rect 253 383 254 384
rect 254 383 255 384
rect 255 383 256 384
rect 256 383 257 384
rect 257 383 258 384
rect 258 383 259 384
rect 259 383 260 384
rect 260 383 261 384
rect 261 383 262 384
rect 262 383 263 384
rect 263 383 264 384
rect 264 383 265 384
rect 265 383 266 384
rect 266 383 267 384
rect 267 383 268 384
rect 268 383 269 384
rect 269 383 270 384
rect 270 383 271 384
rect 271 383 272 384
rect 272 383 273 384
rect 273 383 274 384
rect 274 383 275 384
rect 275 383 276 384
rect 276 383 277 384
rect 277 383 278 384
rect 278 383 279 384
rect 279 383 280 384
rect 280 383 281 384
rect 281 383 282 384
rect 282 383 283 384
rect 283 383 284 384
rect 284 383 285 384
rect 285 383 286 384
rect 286 383 287 384
rect 287 383 288 384
rect 288 383 289 384
rect 289 383 290 384
rect 290 383 291 384
rect 291 383 292 384
rect 292 383 293 384
rect 293 383 294 384
rect 294 383 295 384
rect 295 383 296 384
rect 296 383 297 384
rect 297 383 298 384
rect 298 383 299 384
rect 299 383 300 384
rect 300 383 301 384
rect 301 383 302 384
rect 302 383 303 384
rect 303 383 304 384
rect 304 383 305 384
rect 305 383 306 384
rect 306 383 307 384
rect 307 383 308 384
rect 308 383 309 384
rect 309 383 310 384
rect 310 383 311 384
rect 311 383 312 384
rect 312 383 313 384
rect 313 383 314 384
rect 314 383 315 384
rect 315 383 316 384
rect 316 383 317 384
rect 317 383 318 384
rect 484 383 485 384
rect 485 383 486 384
rect 486 383 487 384
rect 487 383 488 384
rect 488 383 489 384
rect 489 383 490 384
rect 490 383 491 384
rect 491 383 492 384
rect 492 383 493 384
rect 66 382 67 383
rect 67 382 68 383
rect 68 382 69 383
rect 69 382 70 383
rect 70 382 71 383
rect 71 382 72 383
rect 72 382 73 383
rect 73 382 74 383
rect 74 382 75 383
rect 75 382 76 383
rect 202 382 203 383
rect 203 382 204 383
rect 204 382 205 383
rect 205 382 206 383
rect 206 382 207 383
rect 207 382 208 383
rect 208 382 209 383
rect 209 382 210 383
rect 210 382 211 383
rect 211 382 212 383
rect 212 382 213 383
rect 213 382 214 383
rect 214 382 215 383
rect 215 382 216 383
rect 216 382 217 383
rect 217 382 218 383
rect 218 382 219 383
rect 219 382 220 383
rect 220 382 221 383
rect 221 382 222 383
rect 222 382 223 383
rect 223 382 224 383
rect 224 382 225 383
rect 225 382 226 383
rect 226 382 227 383
rect 227 382 228 383
rect 228 382 229 383
rect 229 382 230 383
rect 230 382 231 383
rect 231 382 232 383
rect 232 382 233 383
rect 233 382 234 383
rect 234 382 235 383
rect 235 382 236 383
rect 236 382 237 383
rect 237 382 238 383
rect 238 382 239 383
rect 239 382 240 383
rect 240 382 241 383
rect 241 382 242 383
rect 242 382 243 383
rect 243 382 244 383
rect 244 382 245 383
rect 245 382 246 383
rect 246 382 247 383
rect 247 382 248 383
rect 248 382 249 383
rect 249 382 250 383
rect 250 382 251 383
rect 251 382 252 383
rect 252 382 253 383
rect 253 382 254 383
rect 254 382 255 383
rect 255 382 256 383
rect 256 382 257 383
rect 257 382 258 383
rect 258 382 259 383
rect 259 382 260 383
rect 260 382 261 383
rect 261 382 262 383
rect 262 382 263 383
rect 263 382 264 383
rect 264 382 265 383
rect 265 382 266 383
rect 266 382 267 383
rect 267 382 268 383
rect 268 382 269 383
rect 269 382 270 383
rect 270 382 271 383
rect 271 382 272 383
rect 272 382 273 383
rect 273 382 274 383
rect 274 382 275 383
rect 275 382 276 383
rect 276 382 277 383
rect 277 382 278 383
rect 278 382 279 383
rect 279 382 280 383
rect 280 382 281 383
rect 281 382 282 383
rect 282 382 283 383
rect 283 382 284 383
rect 284 382 285 383
rect 285 382 286 383
rect 286 382 287 383
rect 287 382 288 383
rect 288 382 289 383
rect 289 382 290 383
rect 290 382 291 383
rect 291 382 292 383
rect 292 382 293 383
rect 293 382 294 383
rect 294 382 295 383
rect 295 382 296 383
rect 296 382 297 383
rect 297 382 298 383
rect 298 382 299 383
rect 299 382 300 383
rect 300 382 301 383
rect 301 382 302 383
rect 302 382 303 383
rect 303 382 304 383
rect 304 382 305 383
rect 305 382 306 383
rect 306 382 307 383
rect 307 382 308 383
rect 308 382 309 383
rect 309 382 310 383
rect 310 382 311 383
rect 311 382 312 383
rect 312 382 313 383
rect 313 382 314 383
rect 314 382 315 383
rect 315 382 316 383
rect 316 382 317 383
rect 317 382 318 383
rect 318 382 319 383
rect 484 382 485 383
rect 485 382 486 383
rect 486 382 487 383
rect 487 382 488 383
rect 488 382 489 383
rect 489 382 490 383
rect 490 382 491 383
rect 491 382 492 383
rect 492 382 493 383
rect 65 381 66 382
rect 66 381 67 382
rect 67 381 68 382
rect 68 381 69 382
rect 69 381 70 382
rect 70 381 71 382
rect 71 381 72 382
rect 72 381 73 382
rect 73 381 74 382
rect 74 381 75 382
rect 75 381 76 382
rect 202 381 203 382
rect 203 381 204 382
rect 204 381 205 382
rect 205 381 206 382
rect 206 381 207 382
rect 207 381 208 382
rect 208 381 209 382
rect 209 381 210 382
rect 210 381 211 382
rect 211 381 212 382
rect 212 381 213 382
rect 213 381 214 382
rect 214 381 215 382
rect 215 381 216 382
rect 216 381 217 382
rect 217 381 218 382
rect 218 381 219 382
rect 219 381 220 382
rect 220 381 221 382
rect 221 381 222 382
rect 222 381 223 382
rect 223 381 224 382
rect 224 381 225 382
rect 225 381 226 382
rect 226 381 227 382
rect 227 381 228 382
rect 228 381 229 382
rect 229 381 230 382
rect 230 381 231 382
rect 231 381 232 382
rect 232 381 233 382
rect 233 381 234 382
rect 234 381 235 382
rect 235 381 236 382
rect 236 381 237 382
rect 237 381 238 382
rect 238 381 239 382
rect 239 381 240 382
rect 240 381 241 382
rect 241 381 242 382
rect 242 381 243 382
rect 243 381 244 382
rect 244 381 245 382
rect 245 381 246 382
rect 246 381 247 382
rect 247 381 248 382
rect 248 381 249 382
rect 249 381 250 382
rect 250 381 251 382
rect 251 381 252 382
rect 252 381 253 382
rect 253 381 254 382
rect 254 381 255 382
rect 255 381 256 382
rect 256 381 257 382
rect 257 381 258 382
rect 258 381 259 382
rect 259 381 260 382
rect 260 381 261 382
rect 261 381 262 382
rect 262 381 263 382
rect 263 381 264 382
rect 264 381 265 382
rect 265 381 266 382
rect 266 381 267 382
rect 267 381 268 382
rect 268 381 269 382
rect 269 381 270 382
rect 270 381 271 382
rect 271 381 272 382
rect 272 381 273 382
rect 273 381 274 382
rect 274 381 275 382
rect 275 381 276 382
rect 276 381 277 382
rect 277 381 278 382
rect 278 381 279 382
rect 279 381 280 382
rect 280 381 281 382
rect 281 381 282 382
rect 282 381 283 382
rect 283 381 284 382
rect 284 381 285 382
rect 285 381 286 382
rect 286 381 287 382
rect 287 381 288 382
rect 288 381 289 382
rect 289 381 290 382
rect 290 381 291 382
rect 291 381 292 382
rect 292 381 293 382
rect 293 381 294 382
rect 294 381 295 382
rect 295 381 296 382
rect 296 381 297 382
rect 297 381 298 382
rect 298 381 299 382
rect 299 381 300 382
rect 300 381 301 382
rect 301 381 302 382
rect 302 381 303 382
rect 303 381 304 382
rect 304 381 305 382
rect 305 381 306 382
rect 306 381 307 382
rect 307 381 308 382
rect 308 381 309 382
rect 309 381 310 382
rect 310 381 311 382
rect 311 381 312 382
rect 312 381 313 382
rect 313 381 314 382
rect 314 381 315 382
rect 315 381 316 382
rect 316 381 317 382
rect 317 381 318 382
rect 318 381 319 382
rect 319 381 320 382
rect 320 381 321 382
rect 484 381 485 382
rect 485 381 486 382
rect 486 381 487 382
rect 487 381 488 382
rect 488 381 489 382
rect 489 381 490 382
rect 490 381 491 382
rect 491 381 492 382
rect 492 381 493 382
rect 65 380 66 381
rect 66 380 67 381
rect 67 380 68 381
rect 68 380 69 381
rect 69 380 70 381
rect 70 380 71 381
rect 71 380 72 381
rect 72 380 73 381
rect 73 380 74 381
rect 74 380 75 381
rect 201 380 202 381
rect 202 380 203 381
rect 203 380 204 381
rect 204 380 205 381
rect 205 380 206 381
rect 206 380 207 381
rect 207 380 208 381
rect 208 380 209 381
rect 209 380 210 381
rect 210 380 211 381
rect 211 380 212 381
rect 212 380 213 381
rect 213 380 214 381
rect 214 380 215 381
rect 215 380 216 381
rect 216 380 217 381
rect 217 380 218 381
rect 218 380 219 381
rect 219 380 220 381
rect 220 380 221 381
rect 221 380 222 381
rect 222 380 223 381
rect 223 380 224 381
rect 224 380 225 381
rect 225 380 226 381
rect 226 380 227 381
rect 227 380 228 381
rect 228 380 229 381
rect 229 380 230 381
rect 230 380 231 381
rect 231 380 232 381
rect 232 380 233 381
rect 233 380 234 381
rect 234 380 235 381
rect 235 380 236 381
rect 236 380 237 381
rect 237 380 238 381
rect 238 380 239 381
rect 239 380 240 381
rect 240 380 241 381
rect 241 380 242 381
rect 242 380 243 381
rect 243 380 244 381
rect 244 380 245 381
rect 245 380 246 381
rect 246 380 247 381
rect 247 380 248 381
rect 248 380 249 381
rect 249 380 250 381
rect 250 380 251 381
rect 251 380 252 381
rect 252 380 253 381
rect 253 380 254 381
rect 254 380 255 381
rect 255 380 256 381
rect 256 380 257 381
rect 257 380 258 381
rect 258 380 259 381
rect 259 380 260 381
rect 260 380 261 381
rect 261 380 262 381
rect 262 380 263 381
rect 263 380 264 381
rect 264 380 265 381
rect 265 380 266 381
rect 266 380 267 381
rect 267 380 268 381
rect 268 380 269 381
rect 269 380 270 381
rect 270 380 271 381
rect 271 380 272 381
rect 272 380 273 381
rect 273 380 274 381
rect 274 380 275 381
rect 275 380 276 381
rect 276 380 277 381
rect 277 380 278 381
rect 278 380 279 381
rect 279 380 280 381
rect 280 380 281 381
rect 281 380 282 381
rect 282 380 283 381
rect 283 380 284 381
rect 284 380 285 381
rect 285 380 286 381
rect 286 380 287 381
rect 287 380 288 381
rect 288 380 289 381
rect 289 380 290 381
rect 290 380 291 381
rect 291 380 292 381
rect 292 380 293 381
rect 293 380 294 381
rect 294 380 295 381
rect 295 380 296 381
rect 296 380 297 381
rect 297 380 298 381
rect 298 380 299 381
rect 299 380 300 381
rect 300 380 301 381
rect 301 380 302 381
rect 302 380 303 381
rect 303 380 304 381
rect 304 380 305 381
rect 305 380 306 381
rect 306 380 307 381
rect 307 380 308 381
rect 308 380 309 381
rect 309 380 310 381
rect 310 380 311 381
rect 311 380 312 381
rect 312 380 313 381
rect 313 380 314 381
rect 314 380 315 381
rect 315 380 316 381
rect 316 380 317 381
rect 317 380 318 381
rect 318 380 319 381
rect 319 380 320 381
rect 320 380 321 381
rect 321 380 322 381
rect 484 380 485 381
rect 485 380 486 381
rect 486 380 487 381
rect 487 380 488 381
rect 488 380 489 381
rect 489 380 490 381
rect 490 380 491 381
rect 491 380 492 381
rect 492 380 493 381
rect 64 379 65 380
rect 65 379 66 380
rect 66 379 67 380
rect 67 379 68 380
rect 68 379 69 380
rect 69 379 70 380
rect 70 379 71 380
rect 71 379 72 380
rect 72 379 73 380
rect 73 379 74 380
rect 74 379 75 380
rect 200 379 201 380
rect 201 379 202 380
rect 202 379 203 380
rect 203 379 204 380
rect 204 379 205 380
rect 205 379 206 380
rect 206 379 207 380
rect 207 379 208 380
rect 208 379 209 380
rect 209 379 210 380
rect 210 379 211 380
rect 211 379 212 380
rect 212 379 213 380
rect 213 379 214 380
rect 214 379 215 380
rect 215 379 216 380
rect 216 379 217 380
rect 217 379 218 380
rect 218 379 219 380
rect 219 379 220 380
rect 220 379 221 380
rect 221 379 222 380
rect 222 379 223 380
rect 223 379 224 380
rect 224 379 225 380
rect 225 379 226 380
rect 226 379 227 380
rect 227 379 228 380
rect 228 379 229 380
rect 229 379 230 380
rect 230 379 231 380
rect 231 379 232 380
rect 232 379 233 380
rect 233 379 234 380
rect 234 379 235 380
rect 235 379 236 380
rect 236 379 237 380
rect 237 379 238 380
rect 238 379 239 380
rect 239 379 240 380
rect 240 379 241 380
rect 241 379 242 380
rect 242 379 243 380
rect 243 379 244 380
rect 244 379 245 380
rect 245 379 246 380
rect 246 379 247 380
rect 247 379 248 380
rect 248 379 249 380
rect 249 379 250 380
rect 250 379 251 380
rect 251 379 252 380
rect 252 379 253 380
rect 253 379 254 380
rect 254 379 255 380
rect 255 379 256 380
rect 256 379 257 380
rect 257 379 258 380
rect 258 379 259 380
rect 259 379 260 380
rect 260 379 261 380
rect 261 379 262 380
rect 262 379 263 380
rect 263 379 264 380
rect 264 379 265 380
rect 265 379 266 380
rect 266 379 267 380
rect 267 379 268 380
rect 268 379 269 380
rect 269 379 270 380
rect 270 379 271 380
rect 271 379 272 380
rect 272 379 273 380
rect 273 379 274 380
rect 274 379 275 380
rect 275 379 276 380
rect 276 379 277 380
rect 277 379 278 380
rect 278 379 279 380
rect 279 379 280 380
rect 280 379 281 380
rect 281 379 282 380
rect 282 379 283 380
rect 283 379 284 380
rect 284 379 285 380
rect 285 379 286 380
rect 286 379 287 380
rect 287 379 288 380
rect 288 379 289 380
rect 289 379 290 380
rect 290 379 291 380
rect 291 379 292 380
rect 292 379 293 380
rect 293 379 294 380
rect 294 379 295 380
rect 295 379 296 380
rect 296 379 297 380
rect 297 379 298 380
rect 298 379 299 380
rect 299 379 300 380
rect 300 379 301 380
rect 301 379 302 380
rect 302 379 303 380
rect 303 379 304 380
rect 304 379 305 380
rect 305 379 306 380
rect 306 379 307 380
rect 307 379 308 380
rect 308 379 309 380
rect 309 379 310 380
rect 310 379 311 380
rect 311 379 312 380
rect 312 379 313 380
rect 313 379 314 380
rect 314 379 315 380
rect 315 379 316 380
rect 316 379 317 380
rect 317 379 318 380
rect 318 379 319 380
rect 319 379 320 380
rect 320 379 321 380
rect 321 379 322 380
rect 322 379 323 380
rect 484 379 485 380
rect 485 379 486 380
rect 486 379 487 380
rect 487 379 488 380
rect 488 379 489 380
rect 489 379 490 380
rect 490 379 491 380
rect 491 379 492 380
rect 492 379 493 380
rect 64 378 65 379
rect 65 378 66 379
rect 66 378 67 379
rect 67 378 68 379
rect 68 378 69 379
rect 69 378 70 379
rect 70 378 71 379
rect 71 378 72 379
rect 72 378 73 379
rect 73 378 74 379
rect 199 378 200 379
rect 200 378 201 379
rect 201 378 202 379
rect 202 378 203 379
rect 203 378 204 379
rect 204 378 205 379
rect 205 378 206 379
rect 206 378 207 379
rect 207 378 208 379
rect 208 378 209 379
rect 209 378 210 379
rect 210 378 211 379
rect 211 378 212 379
rect 212 378 213 379
rect 213 378 214 379
rect 214 378 215 379
rect 215 378 216 379
rect 216 378 217 379
rect 217 378 218 379
rect 218 378 219 379
rect 219 378 220 379
rect 220 378 221 379
rect 221 378 222 379
rect 222 378 223 379
rect 223 378 224 379
rect 224 378 225 379
rect 225 378 226 379
rect 226 378 227 379
rect 227 378 228 379
rect 228 378 229 379
rect 229 378 230 379
rect 230 378 231 379
rect 231 378 232 379
rect 232 378 233 379
rect 233 378 234 379
rect 234 378 235 379
rect 235 378 236 379
rect 236 378 237 379
rect 237 378 238 379
rect 238 378 239 379
rect 239 378 240 379
rect 240 378 241 379
rect 241 378 242 379
rect 242 378 243 379
rect 243 378 244 379
rect 244 378 245 379
rect 245 378 246 379
rect 246 378 247 379
rect 247 378 248 379
rect 248 378 249 379
rect 249 378 250 379
rect 250 378 251 379
rect 251 378 252 379
rect 252 378 253 379
rect 253 378 254 379
rect 254 378 255 379
rect 255 378 256 379
rect 256 378 257 379
rect 257 378 258 379
rect 258 378 259 379
rect 259 378 260 379
rect 260 378 261 379
rect 261 378 262 379
rect 262 378 263 379
rect 263 378 264 379
rect 264 378 265 379
rect 265 378 266 379
rect 266 378 267 379
rect 267 378 268 379
rect 268 378 269 379
rect 269 378 270 379
rect 270 378 271 379
rect 271 378 272 379
rect 272 378 273 379
rect 273 378 274 379
rect 274 378 275 379
rect 275 378 276 379
rect 276 378 277 379
rect 277 378 278 379
rect 278 378 279 379
rect 279 378 280 379
rect 280 378 281 379
rect 281 378 282 379
rect 282 378 283 379
rect 283 378 284 379
rect 284 378 285 379
rect 285 378 286 379
rect 286 378 287 379
rect 287 378 288 379
rect 288 378 289 379
rect 289 378 290 379
rect 290 378 291 379
rect 291 378 292 379
rect 292 378 293 379
rect 293 378 294 379
rect 294 378 295 379
rect 295 378 296 379
rect 296 378 297 379
rect 297 378 298 379
rect 298 378 299 379
rect 299 378 300 379
rect 300 378 301 379
rect 301 378 302 379
rect 302 378 303 379
rect 303 378 304 379
rect 304 378 305 379
rect 305 378 306 379
rect 306 378 307 379
rect 307 378 308 379
rect 308 378 309 379
rect 309 378 310 379
rect 310 378 311 379
rect 311 378 312 379
rect 312 378 313 379
rect 313 378 314 379
rect 314 378 315 379
rect 315 378 316 379
rect 316 378 317 379
rect 317 378 318 379
rect 318 378 319 379
rect 319 378 320 379
rect 320 378 321 379
rect 321 378 322 379
rect 322 378 323 379
rect 323 378 324 379
rect 484 378 485 379
rect 485 378 486 379
rect 486 378 487 379
rect 487 378 488 379
rect 488 378 489 379
rect 489 378 490 379
rect 490 378 491 379
rect 491 378 492 379
rect 492 378 493 379
rect 63 377 64 378
rect 64 377 65 378
rect 65 377 66 378
rect 66 377 67 378
rect 67 377 68 378
rect 68 377 69 378
rect 69 377 70 378
rect 70 377 71 378
rect 71 377 72 378
rect 72 377 73 378
rect 199 377 200 378
rect 200 377 201 378
rect 201 377 202 378
rect 202 377 203 378
rect 203 377 204 378
rect 204 377 205 378
rect 205 377 206 378
rect 206 377 207 378
rect 207 377 208 378
rect 208 377 209 378
rect 209 377 210 378
rect 210 377 211 378
rect 211 377 212 378
rect 212 377 213 378
rect 213 377 214 378
rect 214 377 215 378
rect 215 377 216 378
rect 216 377 217 378
rect 217 377 218 378
rect 218 377 219 378
rect 219 377 220 378
rect 220 377 221 378
rect 221 377 222 378
rect 222 377 223 378
rect 223 377 224 378
rect 224 377 225 378
rect 225 377 226 378
rect 226 377 227 378
rect 227 377 228 378
rect 228 377 229 378
rect 229 377 230 378
rect 230 377 231 378
rect 231 377 232 378
rect 232 377 233 378
rect 233 377 234 378
rect 234 377 235 378
rect 235 377 236 378
rect 236 377 237 378
rect 237 377 238 378
rect 238 377 239 378
rect 239 377 240 378
rect 240 377 241 378
rect 241 377 242 378
rect 242 377 243 378
rect 243 377 244 378
rect 244 377 245 378
rect 245 377 246 378
rect 246 377 247 378
rect 247 377 248 378
rect 248 377 249 378
rect 249 377 250 378
rect 250 377 251 378
rect 251 377 252 378
rect 252 377 253 378
rect 253 377 254 378
rect 254 377 255 378
rect 255 377 256 378
rect 256 377 257 378
rect 257 377 258 378
rect 258 377 259 378
rect 259 377 260 378
rect 260 377 261 378
rect 261 377 262 378
rect 262 377 263 378
rect 263 377 264 378
rect 264 377 265 378
rect 265 377 266 378
rect 266 377 267 378
rect 267 377 268 378
rect 268 377 269 378
rect 269 377 270 378
rect 270 377 271 378
rect 271 377 272 378
rect 272 377 273 378
rect 273 377 274 378
rect 274 377 275 378
rect 275 377 276 378
rect 276 377 277 378
rect 277 377 278 378
rect 278 377 279 378
rect 279 377 280 378
rect 280 377 281 378
rect 281 377 282 378
rect 282 377 283 378
rect 283 377 284 378
rect 284 377 285 378
rect 285 377 286 378
rect 286 377 287 378
rect 287 377 288 378
rect 288 377 289 378
rect 289 377 290 378
rect 290 377 291 378
rect 291 377 292 378
rect 292 377 293 378
rect 293 377 294 378
rect 294 377 295 378
rect 295 377 296 378
rect 296 377 297 378
rect 297 377 298 378
rect 298 377 299 378
rect 299 377 300 378
rect 300 377 301 378
rect 301 377 302 378
rect 302 377 303 378
rect 303 377 304 378
rect 304 377 305 378
rect 305 377 306 378
rect 306 377 307 378
rect 307 377 308 378
rect 308 377 309 378
rect 309 377 310 378
rect 310 377 311 378
rect 311 377 312 378
rect 312 377 313 378
rect 313 377 314 378
rect 314 377 315 378
rect 315 377 316 378
rect 316 377 317 378
rect 317 377 318 378
rect 318 377 319 378
rect 319 377 320 378
rect 320 377 321 378
rect 321 377 322 378
rect 322 377 323 378
rect 323 377 324 378
rect 324 377 325 378
rect 325 377 326 378
rect 326 377 327 378
rect 484 377 485 378
rect 485 377 486 378
rect 486 377 487 378
rect 487 377 488 378
rect 488 377 489 378
rect 489 377 490 378
rect 490 377 491 378
rect 491 377 492 378
rect 492 377 493 378
rect 63 376 64 377
rect 64 376 65 377
rect 65 376 66 377
rect 66 376 67 377
rect 67 376 68 377
rect 68 376 69 377
rect 69 376 70 377
rect 70 376 71 377
rect 71 376 72 377
rect 72 376 73 377
rect 198 376 199 377
rect 199 376 200 377
rect 200 376 201 377
rect 201 376 202 377
rect 202 376 203 377
rect 203 376 204 377
rect 204 376 205 377
rect 205 376 206 377
rect 206 376 207 377
rect 207 376 208 377
rect 208 376 209 377
rect 209 376 210 377
rect 210 376 211 377
rect 211 376 212 377
rect 212 376 213 377
rect 213 376 214 377
rect 214 376 215 377
rect 215 376 216 377
rect 216 376 217 377
rect 217 376 218 377
rect 218 376 219 377
rect 219 376 220 377
rect 220 376 221 377
rect 221 376 222 377
rect 222 376 223 377
rect 223 376 224 377
rect 224 376 225 377
rect 225 376 226 377
rect 226 376 227 377
rect 227 376 228 377
rect 228 376 229 377
rect 229 376 230 377
rect 230 376 231 377
rect 231 376 232 377
rect 232 376 233 377
rect 233 376 234 377
rect 234 376 235 377
rect 235 376 236 377
rect 236 376 237 377
rect 237 376 238 377
rect 238 376 239 377
rect 239 376 240 377
rect 240 376 241 377
rect 241 376 242 377
rect 242 376 243 377
rect 243 376 244 377
rect 244 376 245 377
rect 245 376 246 377
rect 246 376 247 377
rect 247 376 248 377
rect 248 376 249 377
rect 249 376 250 377
rect 250 376 251 377
rect 251 376 252 377
rect 252 376 253 377
rect 253 376 254 377
rect 254 376 255 377
rect 255 376 256 377
rect 256 376 257 377
rect 257 376 258 377
rect 258 376 259 377
rect 259 376 260 377
rect 260 376 261 377
rect 261 376 262 377
rect 262 376 263 377
rect 263 376 264 377
rect 264 376 265 377
rect 265 376 266 377
rect 266 376 267 377
rect 267 376 268 377
rect 268 376 269 377
rect 269 376 270 377
rect 270 376 271 377
rect 271 376 272 377
rect 272 376 273 377
rect 273 376 274 377
rect 274 376 275 377
rect 275 376 276 377
rect 276 376 277 377
rect 277 376 278 377
rect 278 376 279 377
rect 279 376 280 377
rect 280 376 281 377
rect 281 376 282 377
rect 282 376 283 377
rect 283 376 284 377
rect 284 376 285 377
rect 285 376 286 377
rect 286 376 287 377
rect 287 376 288 377
rect 288 376 289 377
rect 289 376 290 377
rect 290 376 291 377
rect 291 376 292 377
rect 292 376 293 377
rect 293 376 294 377
rect 294 376 295 377
rect 295 376 296 377
rect 296 376 297 377
rect 297 376 298 377
rect 298 376 299 377
rect 299 376 300 377
rect 300 376 301 377
rect 301 376 302 377
rect 302 376 303 377
rect 303 376 304 377
rect 304 376 305 377
rect 305 376 306 377
rect 306 376 307 377
rect 307 376 308 377
rect 308 376 309 377
rect 309 376 310 377
rect 310 376 311 377
rect 311 376 312 377
rect 312 376 313 377
rect 313 376 314 377
rect 314 376 315 377
rect 315 376 316 377
rect 316 376 317 377
rect 317 376 318 377
rect 318 376 319 377
rect 319 376 320 377
rect 320 376 321 377
rect 321 376 322 377
rect 322 376 323 377
rect 323 376 324 377
rect 324 376 325 377
rect 325 376 326 377
rect 326 376 327 377
rect 327 376 328 377
rect 328 376 329 377
rect 329 376 330 377
rect 484 376 485 377
rect 485 376 486 377
rect 486 376 487 377
rect 487 376 488 377
rect 488 376 489 377
rect 489 376 490 377
rect 490 376 491 377
rect 491 376 492 377
rect 492 376 493 377
rect 62 375 63 376
rect 63 375 64 376
rect 64 375 65 376
rect 65 375 66 376
rect 66 375 67 376
rect 67 375 68 376
rect 68 375 69 376
rect 69 375 70 376
rect 70 375 71 376
rect 71 375 72 376
rect 198 375 199 376
rect 199 375 200 376
rect 200 375 201 376
rect 201 375 202 376
rect 202 375 203 376
rect 203 375 204 376
rect 204 375 205 376
rect 205 375 206 376
rect 206 375 207 376
rect 207 375 208 376
rect 208 375 209 376
rect 209 375 210 376
rect 210 375 211 376
rect 211 375 212 376
rect 212 375 213 376
rect 213 375 214 376
rect 214 375 215 376
rect 215 375 216 376
rect 216 375 217 376
rect 217 375 218 376
rect 218 375 219 376
rect 219 375 220 376
rect 220 375 221 376
rect 221 375 222 376
rect 222 375 223 376
rect 223 375 224 376
rect 224 375 225 376
rect 225 375 226 376
rect 226 375 227 376
rect 227 375 228 376
rect 228 375 229 376
rect 229 375 230 376
rect 230 375 231 376
rect 231 375 232 376
rect 232 375 233 376
rect 233 375 234 376
rect 234 375 235 376
rect 235 375 236 376
rect 236 375 237 376
rect 237 375 238 376
rect 238 375 239 376
rect 239 375 240 376
rect 240 375 241 376
rect 241 375 242 376
rect 242 375 243 376
rect 243 375 244 376
rect 244 375 245 376
rect 245 375 246 376
rect 246 375 247 376
rect 247 375 248 376
rect 248 375 249 376
rect 249 375 250 376
rect 250 375 251 376
rect 251 375 252 376
rect 252 375 253 376
rect 253 375 254 376
rect 254 375 255 376
rect 255 375 256 376
rect 256 375 257 376
rect 257 375 258 376
rect 258 375 259 376
rect 259 375 260 376
rect 260 375 261 376
rect 261 375 262 376
rect 262 375 263 376
rect 263 375 264 376
rect 264 375 265 376
rect 265 375 266 376
rect 266 375 267 376
rect 267 375 268 376
rect 268 375 269 376
rect 269 375 270 376
rect 270 375 271 376
rect 271 375 272 376
rect 272 375 273 376
rect 273 375 274 376
rect 274 375 275 376
rect 275 375 276 376
rect 276 375 277 376
rect 277 375 278 376
rect 278 375 279 376
rect 279 375 280 376
rect 280 375 281 376
rect 281 375 282 376
rect 282 375 283 376
rect 283 375 284 376
rect 284 375 285 376
rect 285 375 286 376
rect 286 375 287 376
rect 287 375 288 376
rect 288 375 289 376
rect 289 375 290 376
rect 290 375 291 376
rect 291 375 292 376
rect 292 375 293 376
rect 307 375 308 376
rect 308 375 309 376
rect 309 375 310 376
rect 310 375 311 376
rect 311 375 312 376
rect 312 375 313 376
rect 313 375 314 376
rect 314 375 315 376
rect 315 375 316 376
rect 316 375 317 376
rect 317 375 318 376
rect 318 375 319 376
rect 319 375 320 376
rect 320 375 321 376
rect 321 375 322 376
rect 322 375 323 376
rect 323 375 324 376
rect 324 375 325 376
rect 325 375 326 376
rect 326 375 327 376
rect 327 375 328 376
rect 328 375 329 376
rect 329 375 330 376
rect 330 375 331 376
rect 331 375 332 376
rect 484 375 485 376
rect 485 375 486 376
rect 486 375 487 376
rect 487 375 488 376
rect 488 375 489 376
rect 489 375 490 376
rect 490 375 491 376
rect 491 375 492 376
rect 492 375 493 376
rect 62 374 63 375
rect 63 374 64 375
rect 64 374 65 375
rect 65 374 66 375
rect 66 374 67 375
rect 67 374 68 375
rect 68 374 69 375
rect 69 374 70 375
rect 70 374 71 375
rect 71 374 72 375
rect 197 374 198 375
rect 198 374 199 375
rect 199 374 200 375
rect 200 374 201 375
rect 201 374 202 375
rect 202 374 203 375
rect 203 374 204 375
rect 204 374 205 375
rect 205 374 206 375
rect 206 374 207 375
rect 207 374 208 375
rect 208 374 209 375
rect 209 374 210 375
rect 210 374 211 375
rect 211 374 212 375
rect 212 374 213 375
rect 213 374 214 375
rect 214 374 215 375
rect 215 374 216 375
rect 216 374 217 375
rect 217 374 218 375
rect 218 374 219 375
rect 219 374 220 375
rect 220 374 221 375
rect 221 374 222 375
rect 222 374 223 375
rect 223 374 224 375
rect 224 374 225 375
rect 225 374 226 375
rect 226 374 227 375
rect 227 374 228 375
rect 228 374 229 375
rect 229 374 230 375
rect 230 374 231 375
rect 231 374 232 375
rect 232 374 233 375
rect 233 374 234 375
rect 234 374 235 375
rect 235 374 236 375
rect 236 374 237 375
rect 237 374 238 375
rect 238 374 239 375
rect 239 374 240 375
rect 240 374 241 375
rect 241 374 242 375
rect 242 374 243 375
rect 243 374 244 375
rect 244 374 245 375
rect 245 374 246 375
rect 246 374 247 375
rect 247 374 248 375
rect 248 374 249 375
rect 249 374 250 375
rect 250 374 251 375
rect 251 374 252 375
rect 252 374 253 375
rect 253 374 254 375
rect 254 374 255 375
rect 255 374 256 375
rect 256 374 257 375
rect 257 374 258 375
rect 258 374 259 375
rect 259 374 260 375
rect 260 374 261 375
rect 261 374 262 375
rect 262 374 263 375
rect 263 374 264 375
rect 264 374 265 375
rect 265 374 266 375
rect 266 374 267 375
rect 267 374 268 375
rect 268 374 269 375
rect 269 374 270 375
rect 270 374 271 375
rect 271 374 272 375
rect 272 374 273 375
rect 273 374 274 375
rect 274 374 275 375
rect 275 374 276 375
rect 276 374 277 375
rect 277 374 278 375
rect 278 374 279 375
rect 279 374 280 375
rect 280 374 281 375
rect 281 374 282 375
rect 282 374 283 375
rect 283 374 284 375
rect 284 374 285 375
rect 285 374 286 375
rect 286 374 287 375
rect 287 374 288 375
rect 288 374 289 375
rect 289 374 290 375
rect 290 374 291 375
rect 311 374 312 375
rect 312 374 313 375
rect 313 374 314 375
rect 314 374 315 375
rect 315 374 316 375
rect 316 374 317 375
rect 317 374 318 375
rect 318 374 319 375
rect 319 374 320 375
rect 320 374 321 375
rect 321 374 322 375
rect 322 374 323 375
rect 323 374 324 375
rect 324 374 325 375
rect 325 374 326 375
rect 326 374 327 375
rect 327 374 328 375
rect 328 374 329 375
rect 329 374 330 375
rect 330 374 331 375
rect 331 374 332 375
rect 332 374 333 375
rect 333 374 334 375
rect 484 374 485 375
rect 485 374 486 375
rect 486 374 487 375
rect 487 374 488 375
rect 488 374 489 375
rect 489 374 490 375
rect 490 374 491 375
rect 491 374 492 375
rect 492 374 493 375
rect 61 373 62 374
rect 62 373 63 374
rect 63 373 64 374
rect 64 373 65 374
rect 65 373 66 374
rect 66 373 67 374
rect 67 373 68 374
rect 68 373 69 374
rect 69 373 70 374
rect 70 373 71 374
rect 197 373 198 374
rect 198 373 199 374
rect 199 373 200 374
rect 200 373 201 374
rect 201 373 202 374
rect 202 373 203 374
rect 203 373 204 374
rect 204 373 205 374
rect 205 373 206 374
rect 206 373 207 374
rect 207 373 208 374
rect 208 373 209 374
rect 209 373 210 374
rect 210 373 211 374
rect 211 373 212 374
rect 212 373 213 374
rect 213 373 214 374
rect 214 373 215 374
rect 215 373 216 374
rect 216 373 217 374
rect 217 373 218 374
rect 218 373 219 374
rect 219 373 220 374
rect 220 373 221 374
rect 221 373 222 374
rect 222 373 223 374
rect 223 373 224 374
rect 224 373 225 374
rect 225 373 226 374
rect 226 373 227 374
rect 227 373 228 374
rect 228 373 229 374
rect 229 373 230 374
rect 230 373 231 374
rect 231 373 232 374
rect 232 373 233 374
rect 233 373 234 374
rect 234 373 235 374
rect 235 373 236 374
rect 236 373 237 374
rect 237 373 238 374
rect 238 373 239 374
rect 239 373 240 374
rect 240 373 241 374
rect 241 373 242 374
rect 242 373 243 374
rect 243 373 244 374
rect 244 373 245 374
rect 245 373 246 374
rect 246 373 247 374
rect 247 373 248 374
rect 248 373 249 374
rect 249 373 250 374
rect 250 373 251 374
rect 251 373 252 374
rect 252 373 253 374
rect 253 373 254 374
rect 254 373 255 374
rect 255 373 256 374
rect 256 373 257 374
rect 257 373 258 374
rect 258 373 259 374
rect 259 373 260 374
rect 260 373 261 374
rect 261 373 262 374
rect 262 373 263 374
rect 263 373 264 374
rect 264 373 265 374
rect 265 373 266 374
rect 266 373 267 374
rect 267 373 268 374
rect 268 373 269 374
rect 269 373 270 374
rect 270 373 271 374
rect 271 373 272 374
rect 272 373 273 374
rect 273 373 274 374
rect 274 373 275 374
rect 275 373 276 374
rect 276 373 277 374
rect 277 373 278 374
rect 278 373 279 374
rect 279 373 280 374
rect 280 373 281 374
rect 281 373 282 374
rect 282 373 283 374
rect 283 373 284 374
rect 284 373 285 374
rect 285 373 286 374
rect 286 373 287 374
rect 287 373 288 374
rect 288 373 289 374
rect 314 373 315 374
rect 315 373 316 374
rect 316 373 317 374
rect 317 373 318 374
rect 318 373 319 374
rect 319 373 320 374
rect 320 373 321 374
rect 321 373 322 374
rect 322 373 323 374
rect 323 373 324 374
rect 324 373 325 374
rect 325 373 326 374
rect 326 373 327 374
rect 327 373 328 374
rect 328 373 329 374
rect 329 373 330 374
rect 330 373 331 374
rect 331 373 332 374
rect 332 373 333 374
rect 333 373 334 374
rect 334 373 335 374
rect 484 373 485 374
rect 485 373 486 374
rect 486 373 487 374
rect 487 373 488 374
rect 488 373 489 374
rect 489 373 490 374
rect 490 373 491 374
rect 491 373 492 374
rect 492 373 493 374
rect 61 372 62 373
rect 62 372 63 373
rect 63 372 64 373
rect 64 372 65 373
rect 65 372 66 373
rect 66 372 67 373
rect 67 372 68 373
rect 68 372 69 373
rect 69 372 70 373
rect 70 372 71 373
rect 196 372 197 373
rect 197 372 198 373
rect 198 372 199 373
rect 199 372 200 373
rect 200 372 201 373
rect 201 372 202 373
rect 202 372 203 373
rect 203 372 204 373
rect 204 372 205 373
rect 205 372 206 373
rect 206 372 207 373
rect 207 372 208 373
rect 208 372 209 373
rect 209 372 210 373
rect 210 372 211 373
rect 211 372 212 373
rect 212 372 213 373
rect 213 372 214 373
rect 214 372 215 373
rect 220 372 221 373
rect 221 372 222 373
rect 222 372 223 373
rect 223 372 224 373
rect 224 372 225 373
rect 225 372 226 373
rect 226 372 227 373
rect 227 372 228 373
rect 228 372 229 373
rect 229 372 230 373
rect 230 372 231 373
rect 231 372 232 373
rect 232 372 233 373
rect 233 372 234 373
rect 234 372 235 373
rect 235 372 236 373
rect 236 372 237 373
rect 237 372 238 373
rect 238 372 239 373
rect 239 372 240 373
rect 240 372 241 373
rect 241 372 242 373
rect 242 372 243 373
rect 243 372 244 373
rect 244 372 245 373
rect 245 372 246 373
rect 246 372 247 373
rect 247 372 248 373
rect 248 372 249 373
rect 249 372 250 373
rect 250 372 251 373
rect 251 372 252 373
rect 252 372 253 373
rect 253 372 254 373
rect 254 372 255 373
rect 255 372 256 373
rect 256 372 257 373
rect 257 372 258 373
rect 258 372 259 373
rect 259 372 260 373
rect 260 372 261 373
rect 261 372 262 373
rect 262 372 263 373
rect 263 372 264 373
rect 264 372 265 373
rect 265 372 266 373
rect 266 372 267 373
rect 267 372 268 373
rect 268 372 269 373
rect 269 372 270 373
rect 270 372 271 373
rect 271 372 272 373
rect 272 372 273 373
rect 273 372 274 373
rect 274 372 275 373
rect 275 372 276 373
rect 276 372 277 373
rect 277 372 278 373
rect 278 372 279 373
rect 279 372 280 373
rect 280 372 281 373
rect 281 372 282 373
rect 282 372 283 373
rect 283 372 284 373
rect 284 372 285 373
rect 285 372 286 373
rect 286 372 287 373
rect 287 372 288 373
rect 317 372 318 373
rect 318 372 319 373
rect 319 372 320 373
rect 320 372 321 373
rect 321 372 322 373
rect 322 372 323 373
rect 323 372 324 373
rect 324 372 325 373
rect 325 372 326 373
rect 326 372 327 373
rect 327 372 328 373
rect 328 372 329 373
rect 329 372 330 373
rect 330 372 331 373
rect 331 372 332 373
rect 332 372 333 373
rect 333 372 334 373
rect 334 372 335 373
rect 335 372 336 373
rect 336 372 337 373
rect 484 372 485 373
rect 485 372 486 373
rect 486 372 487 373
rect 487 372 488 373
rect 488 372 489 373
rect 489 372 490 373
rect 490 372 491 373
rect 491 372 492 373
rect 61 371 62 372
rect 62 371 63 372
rect 63 371 64 372
rect 64 371 65 372
rect 65 371 66 372
rect 66 371 67 372
rect 67 371 68 372
rect 68 371 69 372
rect 69 371 70 372
rect 196 371 197 372
rect 197 371 198 372
rect 198 371 199 372
rect 199 371 200 372
rect 200 371 201 372
rect 201 371 202 372
rect 202 371 203 372
rect 203 371 204 372
rect 204 371 205 372
rect 205 371 206 372
rect 206 371 207 372
rect 207 371 208 372
rect 208 371 209 372
rect 209 371 210 372
rect 210 371 211 372
rect 211 371 212 372
rect 212 371 213 372
rect 221 371 222 372
rect 222 371 223 372
rect 223 371 224 372
rect 224 371 225 372
rect 225 371 226 372
rect 226 371 227 372
rect 227 371 228 372
rect 228 371 229 372
rect 229 371 230 372
rect 230 371 231 372
rect 231 371 232 372
rect 232 371 233 372
rect 233 371 234 372
rect 234 371 235 372
rect 235 371 236 372
rect 236 371 237 372
rect 237 371 238 372
rect 238 371 239 372
rect 239 371 240 372
rect 240 371 241 372
rect 241 371 242 372
rect 242 371 243 372
rect 243 371 244 372
rect 244 371 245 372
rect 245 371 246 372
rect 246 371 247 372
rect 247 371 248 372
rect 248 371 249 372
rect 249 371 250 372
rect 250 371 251 372
rect 251 371 252 372
rect 252 371 253 372
rect 253 371 254 372
rect 254 371 255 372
rect 255 371 256 372
rect 256 371 257 372
rect 257 371 258 372
rect 258 371 259 372
rect 259 371 260 372
rect 260 371 261 372
rect 261 371 262 372
rect 262 371 263 372
rect 263 371 264 372
rect 264 371 265 372
rect 265 371 266 372
rect 266 371 267 372
rect 267 371 268 372
rect 268 371 269 372
rect 269 371 270 372
rect 270 371 271 372
rect 271 371 272 372
rect 272 371 273 372
rect 273 371 274 372
rect 274 371 275 372
rect 277 371 278 372
rect 278 371 279 372
rect 279 371 280 372
rect 280 371 281 372
rect 281 371 282 372
rect 282 371 283 372
rect 283 371 284 372
rect 284 371 285 372
rect 285 371 286 372
rect 286 371 287 372
rect 319 371 320 372
rect 320 371 321 372
rect 321 371 322 372
rect 322 371 323 372
rect 323 371 324 372
rect 324 371 325 372
rect 325 371 326 372
rect 326 371 327 372
rect 327 371 328 372
rect 328 371 329 372
rect 329 371 330 372
rect 330 371 331 372
rect 331 371 332 372
rect 332 371 333 372
rect 333 371 334 372
rect 334 371 335 372
rect 335 371 336 372
rect 336 371 337 372
rect 337 371 338 372
rect 484 371 485 372
rect 485 371 486 372
rect 486 371 487 372
rect 487 371 488 372
rect 488 371 489 372
rect 489 371 490 372
rect 490 371 491 372
rect 491 371 492 372
rect 60 370 61 371
rect 61 370 62 371
rect 62 370 63 371
rect 63 370 64 371
rect 64 370 65 371
rect 65 370 66 371
rect 66 370 67 371
rect 67 370 68 371
rect 68 370 69 371
rect 69 370 70 371
rect 196 370 197 371
rect 197 370 198 371
rect 198 370 199 371
rect 199 370 200 371
rect 200 370 201 371
rect 201 370 202 371
rect 202 370 203 371
rect 203 370 204 371
rect 204 370 205 371
rect 205 370 206 371
rect 206 370 207 371
rect 207 370 208 371
rect 208 370 209 371
rect 209 370 210 371
rect 210 370 211 371
rect 220 370 221 371
rect 221 370 222 371
rect 222 370 223 371
rect 223 370 224 371
rect 224 370 225 371
rect 225 370 226 371
rect 226 370 227 371
rect 227 370 228 371
rect 228 370 229 371
rect 229 370 230 371
rect 230 370 231 371
rect 231 370 232 371
rect 232 370 233 371
rect 233 370 234 371
rect 234 370 235 371
rect 235 370 236 371
rect 236 370 237 371
rect 237 370 238 371
rect 238 370 239 371
rect 239 370 240 371
rect 240 370 241 371
rect 241 370 242 371
rect 242 370 243 371
rect 243 370 244 371
rect 244 370 245 371
rect 245 370 246 371
rect 246 370 247 371
rect 247 370 248 371
rect 248 370 249 371
rect 249 370 250 371
rect 250 370 251 371
rect 251 370 252 371
rect 252 370 253 371
rect 253 370 254 371
rect 254 370 255 371
rect 255 370 256 371
rect 256 370 257 371
rect 257 370 258 371
rect 258 370 259 371
rect 259 370 260 371
rect 260 370 261 371
rect 261 370 262 371
rect 262 370 263 371
rect 263 370 264 371
rect 264 370 265 371
rect 265 370 266 371
rect 266 370 267 371
rect 267 370 268 371
rect 268 370 269 371
rect 269 370 270 371
rect 270 370 271 371
rect 271 370 272 371
rect 272 370 273 371
rect 273 370 274 371
rect 277 370 278 371
rect 278 370 279 371
rect 279 370 280 371
rect 280 370 281 371
rect 281 370 282 371
rect 282 370 283 371
rect 283 370 284 371
rect 284 370 285 371
rect 285 370 286 371
rect 286 370 287 371
rect 321 370 322 371
rect 322 370 323 371
rect 323 370 324 371
rect 324 370 325 371
rect 325 370 326 371
rect 326 370 327 371
rect 327 370 328 371
rect 328 370 329 371
rect 329 370 330 371
rect 330 370 331 371
rect 331 370 332 371
rect 332 370 333 371
rect 333 370 334 371
rect 334 370 335 371
rect 335 370 336 371
rect 336 370 337 371
rect 337 370 338 371
rect 338 370 339 371
rect 483 370 484 371
rect 484 370 485 371
rect 485 370 486 371
rect 486 370 487 371
rect 487 370 488 371
rect 488 370 489 371
rect 489 370 490 371
rect 490 370 491 371
rect 491 370 492 371
rect 60 369 61 370
rect 61 369 62 370
rect 62 369 63 370
rect 63 369 64 370
rect 64 369 65 370
rect 65 369 66 370
rect 66 369 67 370
rect 67 369 68 370
rect 68 369 69 370
rect 196 369 197 370
rect 197 369 198 370
rect 198 369 199 370
rect 199 369 200 370
rect 200 369 201 370
rect 201 369 202 370
rect 202 369 203 370
rect 203 369 204 370
rect 204 369 205 370
rect 205 369 206 370
rect 206 369 207 370
rect 207 369 208 370
rect 208 369 209 370
rect 209 369 210 370
rect 219 369 220 370
rect 220 369 221 370
rect 221 369 222 370
rect 222 369 223 370
rect 223 369 224 370
rect 224 369 225 370
rect 225 369 226 370
rect 226 369 227 370
rect 227 369 228 370
rect 228 369 229 370
rect 229 369 230 370
rect 230 369 231 370
rect 231 369 232 370
rect 232 369 233 370
rect 233 369 234 370
rect 234 369 235 370
rect 235 369 236 370
rect 236 369 237 370
rect 237 369 238 370
rect 238 369 239 370
rect 239 369 240 370
rect 240 369 241 370
rect 241 369 242 370
rect 242 369 243 370
rect 243 369 244 370
rect 244 369 245 370
rect 245 369 246 370
rect 246 369 247 370
rect 247 369 248 370
rect 248 369 249 370
rect 249 369 250 370
rect 250 369 251 370
rect 251 369 252 370
rect 252 369 253 370
rect 253 369 254 370
rect 254 369 255 370
rect 255 369 256 370
rect 256 369 257 370
rect 257 369 258 370
rect 258 369 259 370
rect 259 369 260 370
rect 260 369 261 370
rect 261 369 262 370
rect 262 369 263 370
rect 263 369 264 370
rect 264 369 265 370
rect 265 369 266 370
rect 266 369 267 370
rect 267 369 268 370
rect 268 369 269 370
rect 269 369 270 370
rect 270 369 271 370
rect 271 369 272 370
rect 277 369 278 370
rect 278 369 279 370
rect 279 369 280 370
rect 280 369 281 370
rect 281 369 282 370
rect 282 369 283 370
rect 283 369 284 370
rect 284 369 285 370
rect 285 369 286 370
rect 323 369 324 370
rect 324 369 325 370
rect 325 369 326 370
rect 326 369 327 370
rect 327 369 328 370
rect 328 369 329 370
rect 329 369 330 370
rect 330 369 331 370
rect 331 369 332 370
rect 332 369 333 370
rect 333 369 334 370
rect 334 369 335 370
rect 335 369 336 370
rect 336 369 337 370
rect 337 369 338 370
rect 338 369 339 370
rect 483 369 484 370
rect 484 369 485 370
rect 485 369 486 370
rect 486 369 487 370
rect 487 369 488 370
rect 488 369 489 370
rect 489 369 490 370
rect 490 369 491 370
rect 491 369 492 370
rect 59 368 60 369
rect 60 368 61 369
rect 61 368 62 369
rect 62 368 63 369
rect 63 368 64 369
rect 64 368 65 369
rect 65 368 66 369
rect 66 368 67 369
rect 67 368 68 369
rect 68 368 69 369
rect 195 368 196 369
rect 196 368 197 369
rect 197 368 198 369
rect 198 368 199 369
rect 199 368 200 369
rect 200 368 201 369
rect 201 368 202 369
rect 202 368 203 369
rect 203 368 204 369
rect 204 368 205 369
rect 205 368 206 369
rect 206 368 207 369
rect 207 368 208 369
rect 218 368 219 369
rect 219 368 220 369
rect 220 368 221 369
rect 221 368 222 369
rect 222 368 223 369
rect 223 368 224 369
rect 224 368 225 369
rect 225 368 226 369
rect 226 368 227 369
rect 227 368 228 369
rect 228 368 229 369
rect 229 368 230 369
rect 230 368 231 369
rect 231 368 232 369
rect 232 368 233 369
rect 233 368 234 369
rect 234 368 235 369
rect 235 368 236 369
rect 236 368 237 369
rect 237 368 238 369
rect 238 368 239 369
rect 239 368 240 369
rect 240 368 241 369
rect 241 368 242 369
rect 242 368 243 369
rect 243 368 244 369
rect 244 368 245 369
rect 245 368 246 369
rect 246 368 247 369
rect 247 368 248 369
rect 248 368 249 369
rect 249 368 250 369
rect 250 368 251 369
rect 251 368 252 369
rect 252 368 253 369
rect 253 368 254 369
rect 254 368 255 369
rect 255 368 256 369
rect 256 368 257 369
rect 257 368 258 369
rect 258 368 259 369
rect 259 368 260 369
rect 260 368 261 369
rect 261 368 262 369
rect 262 368 263 369
rect 263 368 264 369
rect 264 368 265 369
rect 265 368 266 369
rect 266 368 267 369
rect 267 368 268 369
rect 268 368 269 369
rect 269 368 270 369
rect 270 368 271 369
rect 277 368 278 369
rect 278 368 279 369
rect 279 368 280 369
rect 280 368 281 369
rect 281 368 282 369
rect 282 368 283 369
rect 283 368 284 369
rect 284 368 285 369
rect 285 368 286 369
rect 324 368 325 369
rect 325 368 326 369
rect 326 368 327 369
rect 327 368 328 369
rect 328 368 329 369
rect 329 368 330 369
rect 330 368 331 369
rect 331 368 332 369
rect 332 368 333 369
rect 333 368 334 369
rect 334 368 335 369
rect 335 368 336 369
rect 336 368 337 369
rect 337 368 338 369
rect 338 368 339 369
rect 339 368 340 369
rect 483 368 484 369
rect 484 368 485 369
rect 485 368 486 369
rect 486 368 487 369
rect 487 368 488 369
rect 488 368 489 369
rect 489 368 490 369
rect 490 368 491 369
rect 491 368 492 369
rect 59 367 60 368
rect 60 367 61 368
rect 61 367 62 368
rect 62 367 63 368
rect 63 367 64 368
rect 64 367 65 368
rect 65 367 66 368
rect 66 367 67 368
rect 67 367 68 368
rect 195 367 196 368
rect 196 367 197 368
rect 197 367 198 368
rect 198 367 199 368
rect 199 367 200 368
rect 200 367 201 368
rect 201 367 202 368
rect 202 367 203 368
rect 203 367 204 368
rect 204 367 205 368
rect 205 367 206 368
rect 206 367 207 368
rect 217 367 218 368
rect 218 367 219 368
rect 219 367 220 368
rect 220 367 221 368
rect 221 367 222 368
rect 222 367 223 368
rect 223 367 224 368
rect 224 367 225 368
rect 225 367 226 368
rect 226 367 227 368
rect 227 367 228 368
rect 228 367 229 368
rect 229 367 230 368
rect 230 367 231 368
rect 231 367 232 368
rect 232 367 233 368
rect 233 367 234 368
rect 234 367 235 368
rect 235 367 236 368
rect 236 367 237 368
rect 237 367 238 368
rect 238 367 239 368
rect 239 367 240 368
rect 240 367 241 368
rect 241 367 242 368
rect 242 367 243 368
rect 243 367 244 368
rect 244 367 245 368
rect 245 367 246 368
rect 246 367 247 368
rect 247 367 248 368
rect 248 367 249 368
rect 249 367 250 368
rect 250 367 251 368
rect 251 367 252 368
rect 252 367 253 368
rect 253 367 254 368
rect 254 367 255 368
rect 255 367 256 368
rect 256 367 257 368
rect 257 367 258 368
rect 258 367 259 368
rect 259 367 260 368
rect 260 367 261 368
rect 261 367 262 368
rect 262 367 263 368
rect 263 367 264 368
rect 264 367 265 368
rect 265 367 266 368
rect 266 367 267 368
rect 267 367 268 368
rect 268 367 269 368
rect 269 367 270 368
rect 277 367 278 368
rect 278 367 279 368
rect 279 367 280 368
rect 280 367 281 368
rect 281 367 282 368
rect 282 367 283 368
rect 283 367 284 368
rect 284 367 285 368
rect 285 367 286 368
rect 326 367 327 368
rect 327 367 328 368
rect 328 367 329 368
rect 329 367 330 368
rect 330 367 331 368
rect 331 367 332 368
rect 332 367 333 368
rect 333 367 334 368
rect 334 367 335 368
rect 335 367 336 368
rect 336 367 337 368
rect 337 367 338 368
rect 338 367 339 368
rect 339 367 340 368
rect 340 367 341 368
rect 483 367 484 368
rect 484 367 485 368
rect 485 367 486 368
rect 486 367 487 368
rect 487 367 488 368
rect 488 367 489 368
rect 489 367 490 368
rect 490 367 491 368
rect 58 366 59 367
rect 59 366 60 367
rect 60 366 61 367
rect 61 366 62 367
rect 62 366 63 367
rect 63 366 64 367
rect 64 366 65 367
rect 65 366 66 367
rect 66 366 67 367
rect 67 366 68 367
rect 195 366 196 367
rect 196 366 197 367
rect 197 366 198 367
rect 198 366 199 367
rect 199 366 200 367
rect 200 366 201 367
rect 201 366 202 367
rect 202 366 203 367
rect 203 366 204 367
rect 204 366 205 367
rect 205 366 206 367
rect 217 366 218 367
rect 218 366 219 367
rect 219 366 220 367
rect 220 366 221 367
rect 221 366 222 367
rect 222 366 223 367
rect 223 366 224 367
rect 224 366 225 367
rect 225 366 226 367
rect 226 366 227 367
rect 227 366 228 367
rect 228 366 229 367
rect 229 366 230 367
rect 230 366 231 367
rect 231 366 232 367
rect 232 366 233 367
rect 233 366 234 367
rect 234 366 235 367
rect 235 366 236 367
rect 236 366 237 367
rect 237 366 238 367
rect 238 366 239 367
rect 239 366 240 367
rect 240 366 241 367
rect 241 366 242 367
rect 242 366 243 367
rect 243 366 244 367
rect 244 366 245 367
rect 245 366 246 367
rect 246 366 247 367
rect 247 366 248 367
rect 248 366 249 367
rect 249 366 250 367
rect 250 366 251 367
rect 251 366 252 367
rect 252 366 253 367
rect 253 366 254 367
rect 254 366 255 367
rect 255 366 256 367
rect 256 366 257 367
rect 257 366 258 367
rect 258 366 259 367
rect 259 366 260 367
rect 260 366 261 367
rect 261 366 262 367
rect 262 366 263 367
rect 263 366 264 367
rect 264 366 265 367
rect 265 366 266 367
rect 266 366 267 367
rect 267 366 268 367
rect 268 366 269 367
rect 278 366 279 367
rect 279 366 280 367
rect 280 366 281 367
rect 281 366 282 367
rect 282 366 283 367
rect 283 366 284 367
rect 284 366 285 367
rect 285 366 286 367
rect 327 366 328 367
rect 328 366 329 367
rect 329 366 330 367
rect 330 366 331 367
rect 331 366 332 367
rect 332 366 333 367
rect 333 366 334 367
rect 334 366 335 367
rect 335 366 336 367
rect 336 366 337 367
rect 337 366 338 367
rect 338 366 339 367
rect 339 366 340 367
rect 340 366 341 367
rect 482 366 483 367
rect 483 366 484 367
rect 484 366 485 367
rect 485 366 486 367
rect 486 366 487 367
rect 487 366 488 367
rect 488 366 489 367
rect 489 366 490 367
rect 490 366 491 367
rect 58 365 59 366
rect 59 365 60 366
rect 60 365 61 366
rect 61 365 62 366
rect 62 365 63 366
rect 63 365 64 366
rect 64 365 65 366
rect 65 365 66 366
rect 66 365 67 366
rect 67 365 68 366
rect 195 365 196 366
rect 196 365 197 366
rect 197 365 198 366
rect 198 365 199 366
rect 199 365 200 366
rect 200 365 201 366
rect 201 365 202 366
rect 202 365 203 366
rect 203 365 204 366
rect 204 365 205 366
rect 205 365 206 366
rect 216 365 217 366
rect 217 365 218 366
rect 218 365 219 366
rect 219 365 220 366
rect 220 365 221 366
rect 221 365 222 366
rect 222 365 223 366
rect 223 365 224 366
rect 224 365 225 366
rect 225 365 226 366
rect 226 365 227 366
rect 227 365 228 366
rect 228 365 229 366
rect 229 365 230 366
rect 230 365 231 366
rect 231 365 232 366
rect 232 365 233 366
rect 233 365 234 366
rect 234 365 235 366
rect 235 365 236 366
rect 236 365 237 366
rect 237 365 238 366
rect 238 365 239 366
rect 239 365 240 366
rect 240 365 241 366
rect 241 365 242 366
rect 242 365 243 366
rect 243 365 244 366
rect 244 365 245 366
rect 245 365 246 366
rect 246 365 247 366
rect 247 365 248 366
rect 248 365 249 366
rect 249 365 250 366
rect 250 365 251 366
rect 251 365 252 366
rect 252 365 253 366
rect 253 365 254 366
rect 254 365 255 366
rect 255 365 256 366
rect 256 365 257 366
rect 257 365 258 366
rect 258 365 259 366
rect 259 365 260 366
rect 260 365 261 366
rect 261 365 262 366
rect 262 365 263 366
rect 263 365 264 366
rect 264 365 265 366
rect 265 365 266 366
rect 266 365 267 366
rect 267 365 268 366
rect 268 365 269 366
rect 278 365 279 366
rect 279 365 280 366
rect 280 365 281 366
rect 281 365 282 366
rect 282 365 283 366
rect 283 365 284 366
rect 284 365 285 366
rect 285 365 286 366
rect 304 365 305 366
rect 305 365 306 366
rect 306 365 307 366
rect 328 365 329 366
rect 329 365 330 366
rect 330 365 331 366
rect 331 365 332 366
rect 332 365 333 366
rect 333 365 334 366
rect 334 365 335 366
rect 335 365 336 366
rect 336 365 337 366
rect 337 365 338 366
rect 338 365 339 366
rect 339 365 340 366
rect 340 365 341 366
rect 341 365 342 366
rect 482 365 483 366
rect 483 365 484 366
rect 484 365 485 366
rect 485 365 486 366
rect 486 365 487 366
rect 487 365 488 366
rect 488 365 489 366
rect 489 365 490 366
rect 490 365 491 366
rect 58 364 59 365
rect 59 364 60 365
rect 60 364 61 365
rect 61 364 62 365
rect 62 364 63 365
rect 63 364 64 365
rect 64 364 65 365
rect 65 364 66 365
rect 66 364 67 365
rect 195 364 196 365
rect 196 364 197 365
rect 197 364 198 365
rect 198 364 199 365
rect 199 364 200 365
rect 200 364 201 365
rect 201 364 202 365
rect 202 364 203 365
rect 203 364 204 365
rect 204 364 205 365
rect 215 364 216 365
rect 216 364 217 365
rect 217 364 218 365
rect 218 364 219 365
rect 219 364 220 365
rect 220 364 221 365
rect 221 364 222 365
rect 222 364 223 365
rect 223 364 224 365
rect 224 364 225 365
rect 225 364 226 365
rect 226 364 227 365
rect 227 364 228 365
rect 228 364 229 365
rect 229 364 230 365
rect 230 364 231 365
rect 231 364 232 365
rect 232 364 233 365
rect 233 364 234 365
rect 234 364 235 365
rect 235 364 236 365
rect 236 364 237 365
rect 237 364 238 365
rect 238 364 239 365
rect 239 364 240 365
rect 240 364 241 365
rect 241 364 242 365
rect 242 364 243 365
rect 246 364 247 365
rect 247 364 248 365
rect 248 364 249 365
rect 249 364 250 365
rect 250 364 251 365
rect 251 364 252 365
rect 252 364 253 365
rect 253 364 254 365
rect 254 364 255 365
rect 255 364 256 365
rect 256 364 257 365
rect 257 364 258 365
rect 258 364 259 365
rect 259 364 260 365
rect 260 364 261 365
rect 261 364 262 365
rect 262 364 263 365
rect 263 364 264 365
rect 264 364 265 365
rect 265 364 266 365
rect 266 364 267 365
rect 267 364 268 365
rect 278 364 279 365
rect 279 364 280 365
rect 280 364 281 365
rect 281 364 282 365
rect 282 364 283 365
rect 283 364 284 365
rect 284 364 285 365
rect 285 364 286 365
rect 300 364 301 365
rect 301 364 302 365
rect 302 364 303 365
rect 303 364 304 365
rect 304 364 305 365
rect 305 364 306 365
rect 306 364 307 365
rect 307 364 308 365
rect 308 364 309 365
rect 309 364 310 365
rect 329 364 330 365
rect 330 364 331 365
rect 331 364 332 365
rect 332 364 333 365
rect 333 364 334 365
rect 334 364 335 365
rect 335 364 336 365
rect 336 364 337 365
rect 337 364 338 365
rect 338 364 339 365
rect 339 364 340 365
rect 340 364 341 365
rect 341 364 342 365
rect 482 364 483 365
rect 483 364 484 365
rect 484 364 485 365
rect 485 364 486 365
rect 486 364 487 365
rect 487 364 488 365
rect 488 364 489 365
rect 489 364 490 365
rect 490 364 491 365
rect 57 363 58 364
rect 58 363 59 364
rect 59 363 60 364
rect 60 363 61 364
rect 61 363 62 364
rect 62 363 63 364
rect 63 363 64 364
rect 64 363 65 364
rect 65 363 66 364
rect 66 363 67 364
rect 195 363 196 364
rect 196 363 197 364
rect 197 363 198 364
rect 198 363 199 364
rect 199 363 200 364
rect 200 363 201 364
rect 201 363 202 364
rect 202 363 203 364
rect 203 363 204 364
rect 214 363 215 364
rect 215 363 216 364
rect 216 363 217 364
rect 217 363 218 364
rect 218 363 219 364
rect 219 363 220 364
rect 220 363 221 364
rect 221 363 222 364
rect 222 363 223 364
rect 223 363 224 364
rect 224 363 225 364
rect 225 363 226 364
rect 226 363 227 364
rect 227 363 228 364
rect 228 363 229 364
rect 229 363 230 364
rect 230 363 231 364
rect 231 363 232 364
rect 232 363 233 364
rect 233 363 234 364
rect 234 363 235 364
rect 235 363 236 364
rect 236 363 237 364
rect 237 363 238 364
rect 238 363 239 364
rect 239 363 240 364
rect 247 363 248 364
rect 248 363 249 364
rect 249 363 250 364
rect 250 363 251 364
rect 251 363 252 364
rect 252 363 253 364
rect 253 363 254 364
rect 254 363 255 364
rect 255 363 256 364
rect 256 363 257 364
rect 257 363 258 364
rect 258 363 259 364
rect 259 363 260 364
rect 260 363 261 364
rect 261 363 262 364
rect 262 363 263 364
rect 263 363 264 364
rect 264 363 265 364
rect 265 363 266 364
rect 266 363 267 364
rect 279 363 280 364
rect 280 363 281 364
rect 281 363 282 364
rect 282 363 283 364
rect 283 363 284 364
rect 284 363 285 364
rect 285 363 286 364
rect 298 363 299 364
rect 299 363 300 364
rect 300 363 301 364
rect 301 363 302 364
rect 302 363 303 364
rect 303 363 304 364
rect 304 363 305 364
rect 305 363 306 364
rect 306 363 307 364
rect 307 363 308 364
rect 308 363 309 364
rect 309 363 310 364
rect 310 363 311 364
rect 311 363 312 364
rect 330 363 331 364
rect 331 363 332 364
rect 332 363 333 364
rect 333 363 334 364
rect 334 363 335 364
rect 335 363 336 364
rect 336 363 337 364
rect 337 363 338 364
rect 338 363 339 364
rect 339 363 340 364
rect 340 363 341 364
rect 341 363 342 364
rect 342 363 343 364
rect 481 363 482 364
rect 482 363 483 364
rect 483 363 484 364
rect 484 363 485 364
rect 485 363 486 364
rect 486 363 487 364
rect 487 363 488 364
rect 488 363 489 364
rect 489 363 490 364
rect 57 362 58 363
rect 58 362 59 363
rect 59 362 60 363
rect 60 362 61 363
rect 61 362 62 363
rect 62 362 63 363
rect 63 362 64 363
rect 64 362 65 363
rect 65 362 66 363
rect 195 362 196 363
rect 196 362 197 363
rect 197 362 198 363
rect 198 362 199 363
rect 199 362 200 363
rect 200 362 201 363
rect 201 362 202 363
rect 202 362 203 363
rect 203 362 204 363
rect 214 362 215 363
rect 215 362 216 363
rect 216 362 217 363
rect 217 362 218 363
rect 218 362 219 363
rect 219 362 220 363
rect 220 362 221 363
rect 221 362 222 363
rect 222 362 223 363
rect 223 362 224 363
rect 224 362 225 363
rect 225 362 226 363
rect 226 362 227 363
rect 227 362 228 363
rect 228 362 229 363
rect 229 362 230 363
rect 230 362 231 363
rect 231 362 232 363
rect 232 362 233 363
rect 233 362 234 363
rect 234 362 235 363
rect 235 362 236 363
rect 236 362 237 363
rect 237 362 238 363
rect 246 362 247 363
rect 247 362 248 363
rect 248 362 249 363
rect 249 362 250 363
rect 250 362 251 363
rect 251 362 252 363
rect 252 362 253 363
rect 253 362 254 363
rect 254 362 255 363
rect 255 362 256 363
rect 256 362 257 363
rect 257 362 258 363
rect 258 362 259 363
rect 259 362 260 363
rect 260 362 261 363
rect 261 362 262 363
rect 262 362 263 363
rect 263 362 264 363
rect 264 362 265 363
rect 265 362 266 363
rect 266 362 267 363
rect 279 362 280 363
rect 280 362 281 363
rect 281 362 282 363
rect 282 362 283 363
rect 283 362 284 363
rect 284 362 285 363
rect 285 362 286 363
rect 286 362 287 363
rect 310 362 311 363
rect 311 362 312 363
rect 312 362 313 363
rect 331 362 332 363
rect 332 362 333 363
rect 333 362 334 363
rect 334 362 335 363
rect 335 362 336 363
rect 336 362 337 363
rect 337 362 338 363
rect 338 362 339 363
rect 339 362 340 363
rect 340 362 341 363
rect 341 362 342 363
rect 342 362 343 363
rect 343 362 344 363
rect 344 362 345 363
rect 345 362 346 363
rect 346 362 347 363
rect 347 362 348 363
rect 481 362 482 363
rect 482 362 483 363
rect 483 362 484 363
rect 484 362 485 363
rect 485 362 486 363
rect 486 362 487 363
rect 487 362 488 363
rect 488 362 489 363
rect 489 362 490 363
rect 57 361 58 362
rect 58 361 59 362
rect 59 361 60 362
rect 60 361 61 362
rect 61 361 62 362
rect 62 361 63 362
rect 63 361 64 362
rect 64 361 65 362
rect 65 361 66 362
rect 195 361 196 362
rect 196 361 197 362
rect 197 361 198 362
rect 198 361 199 362
rect 199 361 200 362
rect 200 361 201 362
rect 201 361 202 362
rect 202 361 203 362
rect 213 361 214 362
rect 214 361 215 362
rect 215 361 216 362
rect 216 361 217 362
rect 217 361 218 362
rect 218 361 219 362
rect 219 361 220 362
rect 220 361 221 362
rect 221 361 222 362
rect 222 361 223 362
rect 223 361 224 362
rect 224 361 225 362
rect 225 361 226 362
rect 226 361 227 362
rect 227 361 228 362
rect 228 361 229 362
rect 229 361 230 362
rect 230 361 231 362
rect 231 361 232 362
rect 232 361 233 362
rect 233 361 234 362
rect 234 361 235 362
rect 235 361 236 362
rect 246 361 247 362
rect 247 361 248 362
rect 248 361 249 362
rect 249 361 250 362
rect 250 361 251 362
rect 251 361 252 362
rect 252 361 253 362
rect 253 361 254 362
rect 254 361 255 362
rect 255 361 256 362
rect 256 361 257 362
rect 257 361 258 362
rect 258 361 259 362
rect 259 361 260 362
rect 260 361 261 362
rect 261 361 262 362
rect 262 361 263 362
rect 263 361 264 362
rect 264 361 265 362
rect 265 361 266 362
rect 280 361 281 362
rect 281 361 282 362
rect 282 361 283 362
rect 283 361 284 362
rect 284 361 285 362
rect 285 361 286 362
rect 286 361 287 362
rect 311 361 312 362
rect 312 361 313 362
rect 313 361 314 362
rect 333 361 334 362
rect 334 361 335 362
rect 335 361 336 362
rect 336 361 337 362
rect 337 361 338 362
rect 338 361 339 362
rect 339 361 340 362
rect 340 361 341 362
rect 341 361 342 362
rect 342 361 343 362
rect 343 361 344 362
rect 344 361 345 362
rect 345 361 346 362
rect 346 361 347 362
rect 347 361 348 362
rect 348 361 349 362
rect 349 361 350 362
rect 350 361 351 362
rect 351 361 352 362
rect 481 361 482 362
rect 482 361 483 362
rect 483 361 484 362
rect 484 361 485 362
rect 485 361 486 362
rect 486 361 487 362
rect 487 361 488 362
rect 488 361 489 362
rect 489 361 490 362
rect 56 360 57 361
rect 57 360 58 361
rect 58 360 59 361
rect 59 360 60 361
rect 60 360 61 361
rect 61 360 62 361
rect 62 360 63 361
rect 63 360 64 361
rect 64 360 65 361
rect 195 360 196 361
rect 196 360 197 361
rect 197 360 198 361
rect 198 360 199 361
rect 199 360 200 361
rect 200 360 201 361
rect 201 360 202 361
rect 202 360 203 361
rect 212 360 213 361
rect 213 360 214 361
rect 214 360 215 361
rect 215 360 216 361
rect 216 360 217 361
rect 217 360 218 361
rect 218 360 219 361
rect 219 360 220 361
rect 220 360 221 361
rect 221 360 222 361
rect 222 360 223 361
rect 223 360 224 361
rect 224 360 225 361
rect 225 360 226 361
rect 226 360 227 361
rect 227 360 228 361
rect 228 360 229 361
rect 229 360 230 361
rect 230 360 231 361
rect 231 360 232 361
rect 232 360 233 361
rect 233 360 234 361
rect 234 360 235 361
rect 245 360 246 361
rect 246 360 247 361
rect 247 360 248 361
rect 248 360 249 361
rect 249 360 250 361
rect 250 360 251 361
rect 251 360 252 361
rect 252 360 253 361
rect 253 360 254 361
rect 254 360 255 361
rect 255 360 256 361
rect 256 360 257 361
rect 257 360 258 361
rect 258 360 259 361
rect 259 360 260 361
rect 260 360 261 361
rect 261 360 262 361
rect 262 360 263 361
rect 263 360 264 361
rect 264 360 265 361
rect 265 360 266 361
rect 280 360 281 361
rect 281 360 282 361
rect 282 360 283 361
rect 283 360 284 361
rect 284 360 285 361
rect 285 360 286 361
rect 286 360 287 361
rect 287 360 288 361
rect 313 360 314 361
rect 314 360 315 361
rect 333 360 334 361
rect 334 360 335 361
rect 335 360 336 361
rect 336 360 337 361
rect 337 360 338 361
rect 338 360 339 361
rect 339 360 340 361
rect 340 360 341 361
rect 341 360 342 361
rect 342 360 343 361
rect 343 360 344 361
rect 344 360 345 361
rect 345 360 346 361
rect 346 360 347 361
rect 347 360 348 361
rect 348 360 349 361
rect 349 360 350 361
rect 350 360 351 361
rect 351 360 352 361
rect 352 360 353 361
rect 353 360 354 361
rect 480 360 481 361
rect 481 360 482 361
rect 482 360 483 361
rect 483 360 484 361
rect 484 360 485 361
rect 485 360 486 361
rect 486 360 487 361
rect 487 360 488 361
rect 488 360 489 361
rect 56 359 57 360
rect 57 359 58 360
rect 58 359 59 360
rect 59 359 60 360
rect 60 359 61 360
rect 61 359 62 360
rect 62 359 63 360
rect 63 359 64 360
rect 64 359 65 360
rect 195 359 196 360
rect 196 359 197 360
rect 197 359 198 360
rect 198 359 199 360
rect 199 359 200 360
rect 200 359 201 360
rect 201 359 202 360
rect 202 359 203 360
rect 212 359 213 360
rect 213 359 214 360
rect 214 359 215 360
rect 215 359 216 360
rect 216 359 217 360
rect 217 359 218 360
rect 218 359 219 360
rect 219 359 220 360
rect 220 359 221 360
rect 221 359 222 360
rect 222 359 223 360
rect 223 359 224 360
rect 224 359 225 360
rect 225 359 226 360
rect 226 359 227 360
rect 227 359 228 360
rect 228 359 229 360
rect 229 359 230 360
rect 230 359 231 360
rect 231 359 232 360
rect 232 359 233 360
rect 233 359 234 360
rect 245 359 246 360
rect 246 359 247 360
rect 247 359 248 360
rect 248 359 249 360
rect 249 359 250 360
rect 250 359 251 360
rect 251 359 252 360
rect 252 359 253 360
rect 253 359 254 360
rect 254 359 255 360
rect 255 359 256 360
rect 256 359 257 360
rect 257 359 258 360
rect 258 359 259 360
rect 259 359 260 360
rect 260 359 261 360
rect 261 359 262 360
rect 262 359 263 360
rect 263 359 264 360
rect 264 359 265 360
rect 281 359 282 360
rect 282 359 283 360
rect 283 359 284 360
rect 284 359 285 360
rect 285 359 286 360
rect 286 359 287 360
rect 287 359 288 360
rect 288 359 289 360
rect 314 359 315 360
rect 334 359 335 360
rect 335 359 336 360
rect 336 359 337 360
rect 337 359 338 360
rect 338 359 339 360
rect 339 359 340 360
rect 340 359 341 360
rect 341 359 342 360
rect 342 359 343 360
rect 343 359 344 360
rect 344 359 345 360
rect 345 359 346 360
rect 346 359 347 360
rect 347 359 348 360
rect 348 359 349 360
rect 349 359 350 360
rect 350 359 351 360
rect 351 359 352 360
rect 352 359 353 360
rect 353 359 354 360
rect 354 359 355 360
rect 355 359 356 360
rect 356 359 357 360
rect 480 359 481 360
rect 481 359 482 360
rect 482 359 483 360
rect 483 359 484 360
rect 484 359 485 360
rect 485 359 486 360
rect 486 359 487 360
rect 487 359 488 360
rect 488 359 489 360
rect 55 358 56 359
rect 56 358 57 359
rect 57 358 58 359
rect 58 358 59 359
rect 59 358 60 359
rect 60 358 61 359
rect 61 358 62 359
rect 62 358 63 359
rect 63 358 64 359
rect 64 358 65 359
rect 194 358 195 359
rect 195 358 196 359
rect 196 358 197 359
rect 197 358 198 359
rect 198 358 199 359
rect 199 358 200 359
rect 200 358 201 359
rect 201 358 202 359
rect 211 358 212 359
rect 212 358 213 359
rect 213 358 214 359
rect 214 358 215 359
rect 215 358 216 359
rect 216 358 217 359
rect 217 358 218 359
rect 218 358 219 359
rect 219 358 220 359
rect 220 358 221 359
rect 221 358 222 359
rect 222 358 223 359
rect 223 358 224 359
rect 224 358 225 359
rect 225 358 226 359
rect 226 358 227 359
rect 227 358 228 359
rect 228 358 229 359
rect 229 358 230 359
rect 230 358 231 359
rect 231 358 232 359
rect 232 358 233 359
rect 244 358 245 359
rect 245 358 246 359
rect 246 358 247 359
rect 247 358 248 359
rect 248 358 249 359
rect 249 358 250 359
rect 250 358 251 359
rect 251 358 252 359
rect 252 358 253 359
rect 253 358 254 359
rect 254 358 255 359
rect 255 358 256 359
rect 256 358 257 359
rect 257 358 258 359
rect 258 358 259 359
rect 259 358 260 359
rect 260 358 261 359
rect 261 358 262 359
rect 262 358 263 359
rect 263 358 264 359
rect 264 358 265 359
rect 282 358 283 359
rect 283 358 284 359
rect 284 358 285 359
rect 285 358 286 359
rect 286 358 287 359
rect 287 358 288 359
rect 288 358 289 359
rect 315 358 316 359
rect 335 358 336 359
rect 336 358 337 359
rect 337 358 338 359
rect 338 358 339 359
rect 339 358 340 359
rect 340 358 341 359
rect 341 358 342 359
rect 342 358 343 359
rect 343 358 344 359
rect 344 358 345 359
rect 345 358 346 359
rect 346 358 347 359
rect 347 358 348 359
rect 348 358 349 359
rect 349 358 350 359
rect 350 358 351 359
rect 351 358 352 359
rect 352 358 353 359
rect 353 358 354 359
rect 354 358 355 359
rect 355 358 356 359
rect 356 358 357 359
rect 357 358 358 359
rect 358 358 359 359
rect 479 358 480 359
rect 480 358 481 359
rect 481 358 482 359
rect 482 358 483 359
rect 483 358 484 359
rect 484 358 485 359
rect 485 358 486 359
rect 486 358 487 359
rect 487 358 488 359
rect 55 357 56 358
rect 56 357 57 358
rect 57 357 58 358
rect 58 357 59 358
rect 59 357 60 358
rect 60 357 61 358
rect 61 357 62 358
rect 62 357 63 358
rect 63 357 64 358
rect 193 357 194 358
rect 194 357 195 358
rect 195 357 196 358
rect 196 357 197 358
rect 197 357 198 358
rect 198 357 199 358
rect 199 357 200 358
rect 200 357 201 358
rect 201 357 202 358
rect 211 357 212 358
rect 212 357 213 358
rect 213 357 214 358
rect 214 357 215 358
rect 215 357 216 358
rect 216 357 217 358
rect 217 357 218 358
rect 218 357 219 358
rect 219 357 220 358
rect 224 357 225 358
rect 225 357 226 358
rect 226 357 227 358
rect 227 357 228 358
rect 228 357 229 358
rect 229 357 230 358
rect 230 357 231 358
rect 231 357 232 358
rect 244 357 245 358
rect 245 357 246 358
rect 246 357 247 358
rect 247 357 248 358
rect 248 357 249 358
rect 249 357 250 358
rect 250 357 251 358
rect 251 357 252 358
rect 252 357 253 358
rect 253 357 254 358
rect 254 357 255 358
rect 255 357 256 358
rect 256 357 257 358
rect 257 357 258 358
rect 258 357 259 358
rect 259 357 260 358
rect 260 357 261 358
rect 261 357 262 358
rect 262 357 263 358
rect 263 357 264 358
rect 283 357 284 358
rect 284 357 285 358
rect 285 357 286 358
rect 286 357 287 358
rect 287 357 288 358
rect 288 357 289 358
rect 289 357 290 358
rect 336 357 337 358
rect 337 357 338 358
rect 338 357 339 358
rect 339 357 340 358
rect 340 357 341 358
rect 341 357 342 358
rect 342 357 343 358
rect 343 357 344 358
rect 344 357 345 358
rect 345 357 346 358
rect 346 357 347 358
rect 347 357 348 358
rect 348 357 349 358
rect 349 357 350 358
rect 350 357 351 358
rect 351 357 352 358
rect 352 357 353 358
rect 353 357 354 358
rect 354 357 355 358
rect 355 357 356 358
rect 356 357 357 358
rect 357 357 358 358
rect 358 357 359 358
rect 359 357 360 358
rect 360 357 361 358
rect 479 357 480 358
rect 480 357 481 358
rect 481 357 482 358
rect 482 357 483 358
rect 483 357 484 358
rect 484 357 485 358
rect 485 357 486 358
rect 486 357 487 358
rect 487 357 488 358
rect 55 356 56 357
rect 56 356 57 357
rect 57 356 58 357
rect 58 356 59 357
rect 59 356 60 357
rect 60 356 61 357
rect 61 356 62 357
rect 62 356 63 357
rect 63 356 64 357
rect 192 356 193 357
rect 193 356 194 357
rect 194 356 195 357
rect 195 356 196 357
rect 196 356 197 357
rect 197 356 198 357
rect 198 356 199 357
rect 199 356 200 357
rect 200 356 201 357
rect 201 356 202 357
rect 210 356 211 357
rect 211 356 212 357
rect 212 356 213 357
rect 213 356 214 357
rect 214 356 215 357
rect 215 356 216 357
rect 216 356 217 357
rect 217 356 218 357
rect 218 356 219 357
rect 224 356 225 357
rect 225 356 226 357
rect 226 356 227 357
rect 227 356 228 357
rect 228 356 229 357
rect 229 356 230 357
rect 230 356 231 357
rect 231 356 232 357
rect 243 356 244 357
rect 244 356 245 357
rect 245 356 246 357
rect 246 356 247 357
rect 247 356 248 357
rect 248 356 249 357
rect 249 356 250 357
rect 250 356 251 357
rect 251 356 252 357
rect 256 356 257 357
rect 257 356 258 357
rect 258 356 259 357
rect 259 356 260 357
rect 260 356 261 357
rect 261 356 262 357
rect 262 356 263 357
rect 284 356 285 357
rect 285 356 286 357
rect 286 356 287 357
rect 287 356 288 357
rect 288 356 289 357
rect 289 356 290 357
rect 290 356 291 357
rect 337 356 338 357
rect 338 356 339 357
rect 339 356 340 357
rect 340 356 341 357
rect 341 356 342 357
rect 342 356 343 357
rect 343 356 344 357
rect 344 356 345 357
rect 345 356 346 357
rect 346 356 347 357
rect 347 356 348 357
rect 348 356 349 357
rect 349 356 350 357
rect 350 356 351 357
rect 351 356 352 357
rect 352 356 353 357
rect 353 356 354 357
rect 354 356 355 357
rect 355 356 356 357
rect 356 356 357 357
rect 357 356 358 357
rect 358 356 359 357
rect 359 356 360 357
rect 360 356 361 357
rect 361 356 362 357
rect 362 356 363 357
rect 479 356 480 357
rect 480 356 481 357
rect 481 356 482 357
rect 482 356 483 357
rect 483 356 484 357
rect 484 356 485 357
rect 485 356 486 357
rect 486 356 487 357
rect 487 356 488 357
rect 55 355 56 356
rect 56 355 57 356
rect 57 355 58 356
rect 58 355 59 356
rect 59 355 60 356
rect 60 355 61 356
rect 61 355 62 356
rect 62 355 63 356
rect 63 355 64 356
rect 190 355 191 356
rect 191 355 192 356
rect 192 355 193 356
rect 193 355 194 356
rect 194 355 195 356
rect 195 355 196 356
rect 196 355 197 356
rect 197 355 198 356
rect 198 355 199 356
rect 199 355 200 356
rect 200 355 201 356
rect 201 355 202 356
rect 210 355 211 356
rect 211 355 212 356
rect 212 355 213 356
rect 213 355 214 356
rect 214 355 215 356
rect 215 355 216 356
rect 216 355 217 356
rect 217 355 218 356
rect 223 355 224 356
rect 224 355 225 356
rect 225 355 226 356
rect 226 355 227 356
rect 227 355 228 356
rect 228 355 229 356
rect 229 355 230 356
rect 230 355 231 356
rect 243 355 244 356
rect 244 355 245 356
rect 245 355 246 356
rect 246 355 247 356
rect 247 355 248 356
rect 248 355 249 356
rect 249 355 250 356
rect 250 355 251 356
rect 257 355 258 356
rect 258 355 259 356
rect 259 355 260 356
rect 260 355 261 356
rect 261 355 262 356
rect 262 355 263 356
rect 286 355 287 356
rect 287 355 288 356
rect 288 355 289 356
rect 289 355 290 356
rect 290 355 291 356
rect 291 355 292 356
rect 338 355 339 356
rect 339 355 340 356
rect 340 355 341 356
rect 341 355 342 356
rect 342 355 343 356
rect 343 355 344 356
rect 344 355 345 356
rect 345 355 346 356
rect 346 355 347 356
rect 347 355 348 356
rect 348 355 349 356
rect 349 355 350 356
rect 350 355 351 356
rect 351 355 352 356
rect 352 355 353 356
rect 353 355 354 356
rect 354 355 355 356
rect 355 355 356 356
rect 356 355 357 356
rect 357 355 358 356
rect 358 355 359 356
rect 359 355 360 356
rect 360 355 361 356
rect 361 355 362 356
rect 362 355 363 356
rect 363 355 364 356
rect 478 355 479 356
rect 479 355 480 356
rect 480 355 481 356
rect 481 355 482 356
rect 482 355 483 356
rect 483 355 484 356
rect 484 355 485 356
rect 485 355 486 356
rect 486 355 487 356
rect 54 354 55 355
rect 55 354 56 355
rect 56 354 57 355
rect 57 354 58 355
rect 58 354 59 355
rect 59 354 60 355
rect 60 354 61 355
rect 61 354 62 355
rect 62 354 63 355
rect 189 354 190 355
rect 190 354 191 355
rect 191 354 192 355
rect 192 354 193 355
rect 193 354 194 355
rect 194 354 195 355
rect 195 354 196 355
rect 197 354 198 355
rect 198 354 199 355
rect 199 354 200 355
rect 200 354 201 355
rect 201 354 202 355
rect 209 354 210 355
rect 210 354 211 355
rect 211 354 212 355
rect 212 354 213 355
rect 213 354 214 355
rect 214 354 215 355
rect 215 354 216 355
rect 216 354 217 355
rect 223 354 224 355
rect 224 354 225 355
rect 225 354 226 355
rect 226 354 227 355
rect 227 354 228 355
rect 228 354 229 355
rect 229 354 230 355
rect 242 354 243 355
rect 243 354 244 355
rect 244 354 245 355
rect 245 354 246 355
rect 246 354 247 355
rect 247 354 248 355
rect 248 354 249 355
rect 249 354 250 355
rect 257 354 258 355
rect 258 354 259 355
rect 259 354 260 355
rect 260 354 261 355
rect 261 354 262 355
rect 338 354 339 355
rect 339 354 340 355
rect 340 354 341 355
rect 341 354 342 355
rect 342 354 343 355
rect 343 354 344 355
rect 344 354 345 355
rect 345 354 346 355
rect 346 354 347 355
rect 347 354 348 355
rect 348 354 349 355
rect 349 354 350 355
rect 350 354 351 355
rect 351 354 352 355
rect 352 354 353 355
rect 353 354 354 355
rect 354 354 355 355
rect 355 354 356 355
rect 356 354 357 355
rect 357 354 358 355
rect 358 354 359 355
rect 359 354 360 355
rect 360 354 361 355
rect 361 354 362 355
rect 362 354 363 355
rect 363 354 364 355
rect 364 354 365 355
rect 478 354 479 355
rect 479 354 480 355
rect 480 354 481 355
rect 481 354 482 355
rect 482 354 483 355
rect 483 354 484 355
rect 484 354 485 355
rect 485 354 486 355
rect 486 354 487 355
rect 54 353 55 354
rect 55 353 56 354
rect 56 353 57 354
rect 57 353 58 354
rect 58 353 59 354
rect 59 353 60 354
rect 60 353 61 354
rect 61 353 62 354
rect 62 353 63 354
rect 188 353 189 354
rect 189 353 190 354
rect 190 353 191 354
rect 191 353 192 354
rect 192 353 193 354
rect 193 353 194 354
rect 194 353 195 354
rect 197 353 198 354
rect 198 353 199 354
rect 199 353 200 354
rect 200 353 201 354
rect 201 353 202 354
rect 209 353 210 354
rect 210 353 211 354
rect 211 353 212 354
rect 212 353 213 354
rect 213 353 214 354
rect 214 353 215 354
rect 215 353 216 354
rect 223 353 224 354
rect 224 353 225 354
rect 225 353 226 354
rect 226 353 227 354
rect 227 353 228 354
rect 228 353 229 354
rect 229 353 230 354
rect 242 353 243 354
rect 243 353 244 354
rect 244 353 245 354
rect 245 353 246 354
rect 246 353 247 354
rect 247 353 248 354
rect 248 353 249 354
rect 256 353 257 354
rect 257 353 258 354
rect 258 353 259 354
rect 259 353 260 354
rect 260 353 261 354
rect 339 353 340 354
rect 340 353 341 354
rect 341 353 342 354
rect 342 353 343 354
rect 343 353 344 354
rect 344 353 345 354
rect 345 353 346 354
rect 346 353 347 354
rect 347 353 348 354
rect 348 353 349 354
rect 349 353 350 354
rect 350 353 351 354
rect 351 353 352 354
rect 352 353 353 354
rect 353 353 354 354
rect 354 353 355 354
rect 355 353 356 354
rect 356 353 357 354
rect 357 353 358 354
rect 358 353 359 354
rect 359 353 360 354
rect 360 353 361 354
rect 361 353 362 354
rect 362 353 363 354
rect 363 353 364 354
rect 364 353 365 354
rect 365 353 366 354
rect 366 353 367 354
rect 477 353 478 354
rect 478 353 479 354
rect 479 353 480 354
rect 480 353 481 354
rect 481 353 482 354
rect 482 353 483 354
rect 483 353 484 354
rect 484 353 485 354
rect 485 353 486 354
rect 54 352 55 353
rect 55 352 56 353
rect 56 352 57 353
rect 57 352 58 353
rect 58 352 59 353
rect 59 352 60 353
rect 60 352 61 353
rect 61 352 62 353
rect 62 352 63 353
rect 188 352 189 353
rect 189 352 190 353
rect 190 352 191 353
rect 191 352 192 353
rect 192 352 193 353
rect 193 352 194 353
rect 198 352 199 353
rect 199 352 200 353
rect 200 352 201 353
rect 201 352 202 353
rect 209 352 210 353
rect 210 352 211 353
rect 211 352 212 353
rect 212 352 213 353
rect 213 352 214 353
rect 214 352 215 353
rect 222 352 223 353
rect 223 352 224 353
rect 224 352 225 353
rect 225 352 226 353
rect 226 352 227 353
rect 227 352 228 353
rect 228 352 229 353
rect 241 352 242 353
rect 242 352 243 353
rect 243 352 244 353
rect 244 352 245 353
rect 245 352 246 353
rect 246 352 247 353
rect 247 352 248 353
rect 255 352 256 353
rect 256 352 257 353
rect 257 352 258 353
rect 258 352 259 353
rect 259 352 260 353
rect 339 352 340 353
rect 340 352 341 353
rect 341 352 342 353
rect 342 352 343 353
rect 343 352 344 353
rect 344 352 345 353
rect 345 352 346 353
rect 346 352 347 353
rect 347 352 348 353
rect 348 352 349 353
rect 349 352 350 353
rect 350 352 351 353
rect 351 352 352 353
rect 352 352 353 353
rect 353 352 354 353
rect 354 352 355 353
rect 355 352 356 353
rect 356 352 357 353
rect 357 352 358 353
rect 358 352 359 353
rect 359 352 360 353
rect 360 352 361 353
rect 361 352 362 353
rect 362 352 363 353
rect 363 352 364 353
rect 364 352 365 353
rect 365 352 366 353
rect 366 352 367 353
rect 367 352 368 353
rect 477 352 478 353
rect 478 352 479 353
rect 479 352 480 353
rect 480 352 481 353
rect 481 352 482 353
rect 482 352 483 353
rect 483 352 484 353
rect 484 352 485 353
rect 485 352 486 353
rect 53 351 54 352
rect 54 351 55 352
rect 55 351 56 352
rect 56 351 57 352
rect 57 351 58 352
rect 58 351 59 352
rect 59 351 60 352
rect 60 351 61 352
rect 61 351 62 352
rect 187 351 188 352
rect 188 351 189 352
rect 189 351 190 352
rect 190 351 191 352
rect 191 351 192 352
rect 192 351 193 352
rect 193 351 194 352
rect 198 351 199 352
rect 199 351 200 352
rect 200 351 201 352
rect 201 351 202 352
rect 209 351 210 352
rect 210 351 211 352
rect 211 351 212 352
rect 212 351 213 352
rect 213 351 214 352
rect 214 351 215 352
rect 222 351 223 352
rect 223 351 224 352
rect 224 351 225 352
rect 225 351 226 352
rect 226 351 227 352
rect 227 351 228 352
rect 241 351 242 352
rect 242 351 243 352
rect 243 351 244 352
rect 244 351 245 352
rect 245 351 246 352
rect 246 351 247 352
rect 254 351 255 352
rect 255 351 256 352
rect 256 351 257 352
rect 257 351 258 352
rect 258 351 259 352
rect 296 351 297 352
rect 297 351 298 352
rect 298 351 299 352
rect 299 351 300 352
rect 300 351 301 352
rect 301 351 302 352
rect 302 351 303 352
rect 340 351 341 352
rect 341 351 342 352
rect 342 351 343 352
rect 343 351 344 352
rect 344 351 345 352
rect 345 351 346 352
rect 346 351 347 352
rect 347 351 348 352
rect 348 351 349 352
rect 349 351 350 352
rect 350 351 351 352
rect 351 351 352 352
rect 352 351 353 352
rect 353 351 354 352
rect 354 351 355 352
rect 355 351 356 352
rect 356 351 357 352
rect 357 351 358 352
rect 358 351 359 352
rect 359 351 360 352
rect 360 351 361 352
rect 361 351 362 352
rect 362 351 363 352
rect 363 351 364 352
rect 364 351 365 352
rect 365 351 366 352
rect 366 351 367 352
rect 367 351 368 352
rect 368 351 369 352
rect 476 351 477 352
rect 477 351 478 352
rect 478 351 479 352
rect 479 351 480 352
rect 480 351 481 352
rect 481 351 482 352
rect 482 351 483 352
rect 483 351 484 352
rect 484 351 485 352
rect 53 350 54 351
rect 54 350 55 351
rect 55 350 56 351
rect 56 350 57 351
rect 57 350 58 351
rect 58 350 59 351
rect 59 350 60 351
rect 60 350 61 351
rect 61 350 62 351
rect 186 350 187 351
rect 187 350 188 351
rect 188 350 189 351
rect 189 350 190 351
rect 190 350 191 351
rect 191 350 192 351
rect 192 350 193 351
rect 199 350 200 351
rect 200 350 201 351
rect 201 350 202 351
rect 209 350 210 351
rect 210 350 211 351
rect 211 350 212 351
rect 212 350 213 351
rect 213 350 214 351
rect 222 350 223 351
rect 223 350 224 351
rect 224 350 225 351
rect 225 350 226 351
rect 226 350 227 351
rect 227 350 228 351
rect 241 350 242 351
rect 242 350 243 351
rect 243 350 244 351
rect 244 350 245 351
rect 245 350 246 351
rect 254 350 255 351
rect 255 350 256 351
rect 256 350 257 351
rect 257 350 258 351
rect 292 350 293 351
rect 293 350 294 351
rect 294 350 295 351
rect 295 350 296 351
rect 296 350 297 351
rect 297 350 298 351
rect 298 350 299 351
rect 299 350 300 351
rect 300 350 301 351
rect 301 350 302 351
rect 302 350 303 351
rect 303 350 304 351
rect 304 350 305 351
rect 305 350 306 351
rect 306 350 307 351
rect 340 350 341 351
rect 341 350 342 351
rect 342 350 343 351
rect 343 350 344 351
rect 344 350 345 351
rect 345 350 346 351
rect 346 350 347 351
rect 347 350 348 351
rect 348 350 349 351
rect 349 350 350 351
rect 350 350 351 351
rect 351 350 352 351
rect 352 350 353 351
rect 353 350 354 351
rect 354 350 355 351
rect 355 350 356 351
rect 356 350 357 351
rect 357 350 358 351
rect 358 350 359 351
rect 359 350 360 351
rect 360 350 361 351
rect 361 350 362 351
rect 362 350 363 351
rect 363 350 364 351
rect 364 350 365 351
rect 365 350 366 351
rect 366 350 367 351
rect 367 350 368 351
rect 368 350 369 351
rect 369 350 370 351
rect 475 350 476 351
rect 476 350 477 351
rect 477 350 478 351
rect 478 350 479 351
rect 479 350 480 351
rect 480 350 481 351
rect 481 350 482 351
rect 482 350 483 351
rect 483 350 484 351
rect 484 350 485 351
rect 53 349 54 350
rect 54 349 55 350
rect 55 349 56 350
rect 56 349 57 350
rect 57 349 58 350
rect 58 349 59 350
rect 59 349 60 350
rect 60 349 61 350
rect 61 349 62 350
rect 186 349 187 350
rect 187 349 188 350
rect 188 349 189 350
rect 189 349 190 350
rect 190 349 191 350
rect 191 349 192 350
rect 199 349 200 350
rect 200 349 201 350
rect 201 349 202 350
rect 209 349 210 350
rect 210 349 211 350
rect 211 349 212 350
rect 212 349 213 350
rect 213 349 214 350
rect 222 349 223 350
rect 223 349 224 350
rect 224 349 225 350
rect 225 349 226 350
rect 226 349 227 350
rect 227 349 228 350
rect 240 349 241 350
rect 241 349 242 350
rect 242 349 243 350
rect 243 349 244 350
rect 244 349 245 350
rect 253 349 254 350
rect 254 349 255 350
rect 255 349 256 350
rect 256 349 257 350
rect 289 349 290 350
rect 290 349 291 350
rect 291 349 292 350
rect 292 349 293 350
rect 293 349 294 350
rect 294 349 295 350
rect 295 349 296 350
rect 296 349 297 350
rect 297 349 298 350
rect 298 349 299 350
rect 299 349 300 350
rect 300 349 301 350
rect 301 349 302 350
rect 302 349 303 350
rect 303 349 304 350
rect 304 349 305 350
rect 305 349 306 350
rect 306 349 307 350
rect 307 349 308 350
rect 308 349 309 350
rect 309 349 310 350
rect 339 349 340 350
rect 340 349 341 350
rect 341 349 342 350
rect 342 349 343 350
rect 343 349 344 350
rect 344 349 345 350
rect 345 349 346 350
rect 346 349 347 350
rect 347 349 348 350
rect 348 349 349 350
rect 349 349 350 350
rect 350 349 351 350
rect 351 349 352 350
rect 352 349 353 350
rect 353 349 354 350
rect 354 349 355 350
rect 355 349 356 350
rect 356 349 357 350
rect 357 349 358 350
rect 358 349 359 350
rect 359 349 360 350
rect 360 349 361 350
rect 361 349 362 350
rect 362 349 363 350
rect 363 349 364 350
rect 364 349 365 350
rect 365 349 366 350
rect 366 349 367 350
rect 367 349 368 350
rect 368 349 369 350
rect 369 349 370 350
rect 475 349 476 350
rect 476 349 477 350
rect 477 349 478 350
rect 478 349 479 350
rect 479 349 480 350
rect 480 349 481 350
rect 481 349 482 350
rect 482 349 483 350
rect 483 349 484 350
rect 52 348 53 349
rect 53 348 54 349
rect 54 348 55 349
rect 55 348 56 349
rect 56 348 57 349
rect 57 348 58 349
rect 58 348 59 349
rect 59 348 60 349
rect 60 348 61 349
rect 186 348 187 349
rect 187 348 188 349
rect 188 348 189 349
rect 189 348 190 349
rect 190 348 191 349
rect 191 348 192 349
rect 200 348 201 349
rect 201 348 202 349
rect 202 348 203 349
rect 209 348 210 349
rect 210 348 211 349
rect 211 348 212 349
rect 212 348 213 349
rect 222 348 223 349
rect 223 348 224 349
rect 224 348 225 349
rect 225 348 226 349
rect 226 348 227 349
rect 240 348 241 349
rect 241 348 242 349
rect 242 348 243 349
rect 243 348 244 349
rect 244 348 245 349
rect 252 348 253 349
rect 253 348 254 349
rect 254 348 255 349
rect 255 348 256 349
rect 288 348 289 349
rect 289 348 290 349
rect 290 348 291 349
rect 291 348 292 349
rect 292 348 293 349
rect 293 348 294 349
rect 294 348 295 349
rect 295 348 296 349
rect 296 348 297 349
rect 303 348 304 349
rect 304 348 305 349
rect 305 348 306 349
rect 306 348 307 349
rect 307 348 308 349
rect 308 348 309 349
rect 309 348 310 349
rect 310 348 311 349
rect 311 348 312 349
rect 339 348 340 349
rect 340 348 341 349
rect 341 348 342 349
rect 342 348 343 349
rect 343 348 344 349
rect 344 348 345 349
rect 345 348 346 349
rect 346 348 347 349
rect 347 348 348 349
rect 348 348 349 349
rect 349 348 350 349
rect 350 348 351 349
rect 351 348 352 349
rect 352 348 353 349
rect 353 348 354 349
rect 354 348 355 349
rect 355 348 356 349
rect 356 348 357 349
rect 357 348 358 349
rect 358 348 359 349
rect 359 348 360 349
rect 360 348 361 349
rect 361 348 362 349
rect 362 348 363 349
rect 363 348 364 349
rect 364 348 365 349
rect 365 348 366 349
rect 366 348 367 349
rect 367 348 368 349
rect 368 348 369 349
rect 369 348 370 349
rect 370 348 371 349
rect 474 348 475 349
rect 475 348 476 349
rect 476 348 477 349
rect 477 348 478 349
rect 478 348 479 349
rect 479 348 480 349
rect 480 348 481 349
rect 481 348 482 349
rect 482 348 483 349
rect 483 348 484 349
rect 52 347 53 348
rect 53 347 54 348
rect 54 347 55 348
rect 55 347 56 348
rect 56 347 57 348
rect 57 347 58 348
rect 58 347 59 348
rect 59 347 60 348
rect 60 347 61 348
rect 185 347 186 348
rect 186 347 187 348
rect 187 347 188 348
rect 188 347 189 348
rect 189 347 190 348
rect 190 347 191 348
rect 191 347 192 348
rect 201 347 202 348
rect 202 347 203 348
rect 209 347 210 348
rect 210 347 211 348
rect 211 347 212 348
rect 212 347 213 348
rect 222 347 223 348
rect 223 347 224 348
rect 224 347 225 348
rect 225 347 226 348
rect 226 347 227 348
rect 240 347 241 348
rect 241 347 242 348
rect 242 347 243 348
rect 243 347 244 348
rect 251 347 252 348
rect 252 347 253 348
rect 253 347 254 348
rect 286 347 287 348
rect 287 347 288 348
rect 288 347 289 348
rect 289 347 290 348
rect 290 347 291 348
rect 308 347 309 348
rect 309 347 310 348
rect 310 347 311 348
rect 311 347 312 348
rect 312 347 313 348
rect 313 347 314 348
rect 339 347 340 348
rect 340 347 341 348
rect 341 347 342 348
rect 342 347 343 348
rect 343 347 344 348
rect 344 347 345 348
rect 345 347 346 348
rect 346 347 347 348
rect 347 347 348 348
rect 348 347 349 348
rect 349 347 350 348
rect 350 347 351 348
rect 351 347 352 348
rect 352 347 353 348
rect 353 347 354 348
rect 354 347 355 348
rect 355 347 356 348
rect 356 347 357 348
rect 357 347 358 348
rect 358 347 359 348
rect 359 347 360 348
rect 360 347 361 348
rect 361 347 362 348
rect 362 347 363 348
rect 363 347 364 348
rect 364 347 365 348
rect 365 347 366 348
rect 366 347 367 348
rect 367 347 368 348
rect 368 347 369 348
rect 369 347 370 348
rect 370 347 371 348
rect 371 347 372 348
rect 474 347 475 348
rect 475 347 476 348
rect 476 347 477 348
rect 477 347 478 348
rect 478 347 479 348
rect 479 347 480 348
rect 480 347 481 348
rect 481 347 482 348
rect 482 347 483 348
rect 52 346 53 347
rect 53 346 54 347
rect 54 346 55 347
rect 55 346 56 347
rect 56 346 57 347
rect 57 346 58 347
rect 58 346 59 347
rect 59 346 60 347
rect 60 346 61 347
rect 183 346 184 347
rect 184 346 185 347
rect 185 346 186 347
rect 186 346 187 347
rect 187 346 188 347
rect 188 346 189 347
rect 189 346 190 347
rect 190 346 191 347
rect 191 346 192 347
rect 202 346 203 347
rect 209 346 210 347
rect 210 346 211 347
rect 211 346 212 347
rect 212 346 213 347
rect 222 346 223 347
rect 223 346 224 347
rect 224 346 225 347
rect 225 346 226 347
rect 240 346 241 347
rect 241 346 242 347
rect 242 346 243 347
rect 250 346 251 347
rect 251 346 252 347
rect 285 346 286 347
rect 286 346 287 347
rect 287 346 288 347
rect 288 346 289 347
rect 311 346 312 347
rect 312 346 313 347
rect 313 346 314 347
rect 314 346 315 347
rect 338 346 339 347
rect 339 346 340 347
rect 340 346 341 347
rect 341 346 342 347
rect 342 346 343 347
rect 343 346 344 347
rect 344 346 345 347
rect 345 346 346 347
rect 346 346 347 347
rect 347 346 348 347
rect 348 346 349 347
rect 349 346 350 347
rect 350 346 351 347
rect 351 346 352 347
rect 352 346 353 347
rect 353 346 354 347
rect 354 346 355 347
rect 355 346 356 347
rect 356 346 357 347
rect 357 346 358 347
rect 358 346 359 347
rect 359 346 360 347
rect 360 346 361 347
rect 361 346 362 347
rect 362 346 363 347
rect 363 346 364 347
rect 364 346 365 347
rect 365 346 366 347
rect 366 346 367 347
rect 367 346 368 347
rect 368 346 369 347
rect 369 346 370 347
rect 370 346 371 347
rect 371 346 372 347
rect 473 346 474 347
rect 474 346 475 347
rect 475 346 476 347
rect 476 346 477 347
rect 477 346 478 347
rect 478 346 479 347
rect 479 346 480 347
rect 480 346 481 347
rect 481 346 482 347
rect 52 345 53 346
rect 53 345 54 346
rect 54 345 55 346
rect 55 345 56 346
rect 56 345 57 346
rect 57 345 58 346
rect 58 345 59 346
rect 59 345 60 346
rect 60 345 61 346
rect 181 345 182 346
rect 182 345 183 346
rect 183 345 184 346
rect 184 345 185 346
rect 185 345 186 346
rect 186 345 187 346
rect 187 345 188 346
rect 188 345 189 346
rect 189 345 190 346
rect 190 345 191 346
rect 191 345 192 346
rect 209 345 210 346
rect 210 345 211 346
rect 211 345 212 346
rect 222 345 223 346
rect 223 345 224 346
rect 224 345 225 346
rect 225 345 226 346
rect 239 345 240 346
rect 240 345 241 346
rect 241 345 242 346
rect 242 345 243 346
rect 249 345 250 346
rect 284 345 285 346
rect 285 345 286 346
rect 286 345 287 346
rect 313 345 314 346
rect 314 345 315 346
rect 315 345 316 346
rect 337 345 338 346
rect 338 345 339 346
rect 339 345 340 346
rect 340 345 341 346
rect 341 345 342 346
rect 342 345 343 346
rect 343 345 344 346
rect 344 345 345 346
rect 345 345 346 346
rect 346 345 347 346
rect 347 345 348 346
rect 348 345 349 346
rect 349 345 350 346
rect 350 345 351 346
rect 351 345 352 346
rect 352 345 353 346
rect 353 345 354 346
rect 354 345 355 346
rect 355 345 356 346
rect 356 345 357 346
rect 357 345 358 346
rect 358 345 359 346
rect 359 345 360 346
rect 360 345 361 346
rect 361 345 362 346
rect 362 345 363 346
rect 363 345 364 346
rect 364 345 365 346
rect 365 345 366 346
rect 366 345 367 346
rect 367 345 368 346
rect 368 345 369 346
rect 369 345 370 346
rect 370 345 371 346
rect 371 345 372 346
rect 372 345 373 346
rect 472 345 473 346
rect 473 345 474 346
rect 474 345 475 346
rect 475 345 476 346
rect 476 345 477 346
rect 477 345 478 346
rect 478 345 479 346
rect 479 345 480 346
rect 480 345 481 346
rect 481 345 482 346
rect 51 344 52 345
rect 52 344 53 345
rect 53 344 54 345
rect 54 344 55 345
rect 55 344 56 345
rect 56 344 57 345
rect 57 344 58 345
rect 58 344 59 345
rect 59 344 60 345
rect 180 344 181 345
rect 181 344 182 345
rect 182 344 183 345
rect 183 344 184 345
rect 184 344 185 345
rect 185 344 186 345
rect 186 344 187 345
rect 187 344 188 345
rect 188 344 189 345
rect 189 344 190 345
rect 190 344 191 345
rect 191 344 192 345
rect 192 344 193 345
rect 210 344 211 345
rect 211 344 212 345
rect 222 344 223 345
rect 223 344 224 345
rect 224 344 225 345
rect 225 344 226 345
rect 239 344 240 345
rect 240 344 241 345
rect 241 344 242 345
rect 283 344 284 345
rect 284 344 285 345
rect 315 344 316 345
rect 316 344 317 345
rect 317 344 318 345
rect 337 344 338 345
rect 338 344 339 345
rect 339 344 340 345
rect 340 344 341 345
rect 341 344 342 345
rect 342 344 343 345
rect 343 344 344 345
rect 344 344 345 345
rect 345 344 346 345
rect 346 344 347 345
rect 347 344 348 345
rect 348 344 349 345
rect 349 344 350 345
rect 350 344 351 345
rect 351 344 352 345
rect 352 344 353 345
rect 353 344 354 345
rect 354 344 355 345
rect 355 344 356 345
rect 356 344 357 345
rect 357 344 358 345
rect 358 344 359 345
rect 359 344 360 345
rect 360 344 361 345
rect 361 344 362 345
rect 362 344 363 345
rect 363 344 364 345
rect 364 344 365 345
rect 365 344 366 345
rect 366 344 367 345
rect 367 344 368 345
rect 368 344 369 345
rect 369 344 370 345
rect 370 344 371 345
rect 371 344 372 345
rect 372 344 373 345
rect 472 344 473 345
rect 473 344 474 345
rect 474 344 475 345
rect 475 344 476 345
rect 476 344 477 345
rect 477 344 478 345
rect 478 344 479 345
rect 479 344 480 345
rect 480 344 481 345
rect 51 343 52 344
rect 52 343 53 344
rect 53 343 54 344
rect 54 343 55 344
rect 55 343 56 344
rect 56 343 57 344
rect 57 343 58 344
rect 58 343 59 344
rect 59 343 60 344
rect 179 343 180 344
rect 180 343 181 344
rect 181 343 182 344
rect 182 343 183 344
rect 183 343 184 344
rect 184 343 185 344
rect 185 343 186 344
rect 186 343 187 344
rect 187 343 188 344
rect 188 343 189 344
rect 189 343 190 344
rect 190 343 191 344
rect 191 343 192 344
rect 192 343 193 344
rect 193 343 194 344
rect 210 343 211 344
rect 211 343 212 344
rect 222 343 223 344
rect 223 343 224 344
rect 224 343 225 344
rect 239 343 240 344
rect 240 343 241 344
rect 241 343 242 344
rect 283 343 284 344
rect 316 343 317 344
rect 317 343 318 344
rect 318 343 319 344
rect 336 343 337 344
rect 337 343 338 344
rect 338 343 339 344
rect 339 343 340 344
rect 340 343 341 344
rect 341 343 342 344
rect 342 343 343 344
rect 343 343 344 344
rect 344 343 345 344
rect 345 343 346 344
rect 346 343 347 344
rect 347 343 348 344
rect 348 343 349 344
rect 349 343 350 344
rect 350 343 351 344
rect 351 343 352 344
rect 352 343 353 344
rect 353 343 354 344
rect 354 343 355 344
rect 355 343 356 344
rect 356 343 357 344
rect 357 343 358 344
rect 358 343 359 344
rect 359 343 360 344
rect 360 343 361 344
rect 361 343 362 344
rect 362 343 363 344
rect 363 343 364 344
rect 364 343 365 344
rect 365 343 366 344
rect 366 343 367 344
rect 367 343 368 344
rect 368 343 369 344
rect 369 343 370 344
rect 370 343 371 344
rect 371 343 372 344
rect 372 343 373 344
rect 373 343 374 344
rect 471 343 472 344
rect 472 343 473 344
rect 473 343 474 344
rect 474 343 475 344
rect 475 343 476 344
rect 476 343 477 344
rect 477 343 478 344
rect 478 343 479 344
rect 479 343 480 344
rect 51 342 52 343
rect 52 342 53 343
rect 53 342 54 343
rect 54 342 55 343
rect 55 342 56 343
rect 56 342 57 343
rect 57 342 58 343
rect 58 342 59 343
rect 59 342 60 343
rect 179 342 180 343
rect 180 342 181 343
rect 181 342 182 343
rect 182 342 183 343
rect 183 342 184 343
rect 184 342 185 343
rect 185 342 186 343
rect 189 342 190 343
rect 190 342 191 343
rect 191 342 192 343
rect 192 342 193 343
rect 193 342 194 343
rect 194 342 195 343
rect 211 342 212 343
rect 222 342 223 343
rect 223 342 224 343
rect 224 342 225 343
rect 239 342 240 343
rect 240 342 241 343
rect 318 342 319 343
rect 319 342 320 343
rect 335 342 336 343
rect 336 342 337 343
rect 337 342 338 343
rect 338 342 339 343
rect 339 342 340 343
rect 340 342 341 343
rect 341 342 342 343
rect 342 342 343 343
rect 343 342 344 343
rect 344 342 345 343
rect 345 342 346 343
rect 346 342 347 343
rect 347 342 348 343
rect 348 342 349 343
rect 349 342 350 343
rect 350 342 351 343
rect 351 342 352 343
rect 352 342 353 343
rect 353 342 354 343
rect 354 342 355 343
rect 355 342 356 343
rect 356 342 357 343
rect 357 342 358 343
rect 358 342 359 343
rect 359 342 360 343
rect 360 342 361 343
rect 361 342 362 343
rect 362 342 363 343
rect 363 342 364 343
rect 364 342 365 343
rect 365 342 366 343
rect 366 342 367 343
rect 367 342 368 343
rect 368 342 369 343
rect 369 342 370 343
rect 370 342 371 343
rect 371 342 372 343
rect 372 342 373 343
rect 373 342 374 343
rect 470 342 471 343
rect 471 342 472 343
rect 472 342 473 343
rect 473 342 474 343
rect 474 342 475 343
rect 475 342 476 343
rect 476 342 477 343
rect 477 342 478 343
rect 478 342 479 343
rect 479 342 480 343
rect 51 341 52 342
rect 52 341 53 342
rect 53 341 54 342
rect 54 341 55 342
rect 55 341 56 342
rect 56 341 57 342
rect 57 341 58 342
rect 58 341 59 342
rect 59 341 60 342
rect 178 341 179 342
rect 179 341 180 342
rect 180 341 181 342
rect 181 341 182 342
rect 182 341 183 342
rect 183 341 184 342
rect 184 341 185 342
rect 190 341 191 342
rect 191 341 192 342
rect 192 341 193 342
rect 193 341 194 342
rect 194 341 195 342
rect 195 341 196 342
rect 223 341 224 342
rect 224 341 225 342
rect 239 341 240 342
rect 240 341 241 342
rect 302 341 303 342
rect 303 341 304 342
rect 319 341 320 342
rect 334 341 335 342
rect 335 341 336 342
rect 336 341 337 342
rect 337 341 338 342
rect 338 341 339 342
rect 339 341 340 342
rect 340 341 341 342
rect 341 341 342 342
rect 342 341 343 342
rect 343 341 344 342
rect 344 341 345 342
rect 345 341 346 342
rect 346 341 347 342
rect 347 341 348 342
rect 348 341 349 342
rect 349 341 350 342
rect 350 341 351 342
rect 351 341 352 342
rect 352 341 353 342
rect 353 341 354 342
rect 354 341 355 342
rect 355 341 356 342
rect 356 341 357 342
rect 357 341 358 342
rect 358 341 359 342
rect 359 341 360 342
rect 360 341 361 342
rect 361 341 362 342
rect 362 341 363 342
rect 363 341 364 342
rect 364 341 365 342
rect 365 341 366 342
rect 366 341 367 342
rect 367 341 368 342
rect 368 341 369 342
rect 369 341 370 342
rect 370 341 371 342
rect 371 341 372 342
rect 372 341 373 342
rect 373 341 374 342
rect 469 341 470 342
rect 470 341 471 342
rect 471 341 472 342
rect 472 341 473 342
rect 473 341 474 342
rect 474 341 475 342
rect 475 341 476 342
rect 476 341 477 342
rect 477 341 478 342
rect 478 341 479 342
rect 50 340 51 341
rect 51 340 52 341
rect 52 340 53 341
rect 53 340 54 341
rect 54 340 55 341
rect 55 340 56 341
rect 56 340 57 341
rect 57 340 58 341
rect 58 340 59 341
rect 178 340 179 341
rect 179 340 180 341
rect 180 340 181 341
rect 181 340 182 341
rect 182 340 183 341
rect 183 340 184 341
rect 191 340 192 341
rect 192 340 193 341
rect 193 340 194 341
rect 194 340 195 341
rect 195 340 196 341
rect 196 340 197 341
rect 223 340 224 341
rect 224 340 225 341
rect 239 340 240 341
rect 302 340 303 341
rect 303 340 304 341
rect 320 340 321 341
rect 333 340 334 341
rect 334 340 335 341
rect 335 340 336 341
rect 336 340 337 341
rect 337 340 338 341
rect 338 340 339 341
rect 339 340 340 341
rect 341 340 342 341
rect 342 340 343 341
rect 343 340 344 341
rect 344 340 345 341
rect 345 340 346 341
rect 346 340 347 341
rect 347 340 348 341
rect 348 340 349 341
rect 349 340 350 341
rect 350 340 351 341
rect 351 340 352 341
rect 352 340 353 341
rect 353 340 354 341
rect 354 340 355 341
rect 355 340 356 341
rect 356 340 357 341
rect 357 340 358 341
rect 358 340 359 341
rect 359 340 360 341
rect 360 340 361 341
rect 361 340 362 341
rect 362 340 363 341
rect 363 340 364 341
rect 364 340 365 341
rect 365 340 366 341
rect 366 340 367 341
rect 367 340 368 341
rect 368 340 369 341
rect 369 340 370 341
rect 370 340 371 341
rect 371 340 372 341
rect 372 340 373 341
rect 373 340 374 341
rect 374 340 375 341
rect 469 340 470 341
rect 470 340 471 341
rect 471 340 472 341
rect 472 340 473 341
rect 473 340 474 341
rect 474 340 475 341
rect 475 340 476 341
rect 476 340 477 341
rect 477 340 478 341
rect 50 339 51 340
rect 51 339 52 340
rect 52 339 53 340
rect 53 339 54 340
rect 54 339 55 340
rect 55 339 56 340
rect 56 339 57 340
rect 57 339 58 340
rect 58 339 59 340
rect 168 339 169 340
rect 177 339 178 340
rect 178 339 179 340
rect 179 339 180 340
rect 180 339 181 340
rect 181 339 182 340
rect 182 339 183 340
rect 193 339 194 340
rect 194 339 195 340
rect 195 339 196 340
rect 196 339 197 340
rect 197 339 198 340
rect 301 339 302 340
rect 302 339 303 340
rect 303 339 304 340
rect 333 339 334 340
rect 334 339 335 340
rect 335 339 336 340
rect 336 339 337 340
rect 337 339 338 340
rect 340 339 341 340
rect 341 339 342 340
rect 342 339 343 340
rect 343 339 344 340
rect 344 339 345 340
rect 345 339 346 340
rect 346 339 347 340
rect 347 339 348 340
rect 348 339 349 340
rect 349 339 350 340
rect 350 339 351 340
rect 351 339 352 340
rect 352 339 353 340
rect 353 339 354 340
rect 354 339 355 340
rect 355 339 356 340
rect 356 339 357 340
rect 357 339 358 340
rect 358 339 359 340
rect 359 339 360 340
rect 360 339 361 340
rect 361 339 362 340
rect 362 339 363 340
rect 363 339 364 340
rect 364 339 365 340
rect 365 339 366 340
rect 366 339 367 340
rect 367 339 368 340
rect 368 339 369 340
rect 369 339 370 340
rect 370 339 371 340
rect 371 339 372 340
rect 372 339 373 340
rect 373 339 374 340
rect 374 339 375 340
rect 468 339 469 340
rect 469 339 470 340
rect 470 339 471 340
rect 471 339 472 340
rect 472 339 473 340
rect 473 339 474 340
rect 474 339 475 340
rect 475 339 476 340
rect 476 339 477 340
rect 477 339 478 340
rect 50 338 51 339
rect 51 338 52 339
rect 52 338 53 339
rect 53 338 54 339
rect 54 338 55 339
rect 55 338 56 339
rect 56 338 57 339
rect 57 338 58 339
rect 58 338 59 339
rect 161 338 162 339
rect 168 338 169 339
rect 169 338 170 339
rect 177 338 178 339
rect 178 338 179 339
rect 179 338 180 339
rect 180 338 181 339
rect 181 338 182 339
rect 182 338 183 339
rect 194 338 195 339
rect 195 338 196 339
rect 196 338 197 339
rect 197 338 198 339
rect 198 338 199 339
rect 288 338 289 339
rect 289 338 290 339
rect 300 338 301 339
rect 301 338 302 339
rect 302 338 303 339
rect 303 338 304 339
rect 332 338 333 339
rect 333 338 334 339
rect 334 338 335 339
rect 335 338 336 339
rect 340 338 341 339
rect 341 338 342 339
rect 342 338 343 339
rect 343 338 344 339
rect 344 338 345 339
rect 345 338 346 339
rect 346 338 347 339
rect 347 338 348 339
rect 348 338 349 339
rect 349 338 350 339
rect 350 338 351 339
rect 351 338 352 339
rect 352 338 353 339
rect 353 338 354 339
rect 354 338 355 339
rect 355 338 356 339
rect 356 338 357 339
rect 357 338 358 339
rect 358 338 359 339
rect 359 338 360 339
rect 360 338 361 339
rect 361 338 362 339
rect 362 338 363 339
rect 363 338 364 339
rect 364 338 365 339
rect 365 338 366 339
rect 366 338 367 339
rect 367 338 368 339
rect 368 338 369 339
rect 369 338 370 339
rect 370 338 371 339
rect 371 338 372 339
rect 372 338 373 339
rect 373 338 374 339
rect 374 338 375 339
rect 467 338 468 339
rect 468 338 469 339
rect 469 338 470 339
rect 470 338 471 339
rect 471 338 472 339
rect 472 338 473 339
rect 473 338 474 339
rect 474 338 475 339
rect 475 338 476 339
rect 476 338 477 339
rect 50 337 51 338
rect 51 337 52 338
rect 52 337 53 338
rect 53 337 54 338
rect 54 337 55 338
rect 55 337 56 338
rect 56 337 57 338
rect 57 337 58 338
rect 58 337 59 338
rect 161 337 162 338
rect 168 337 169 338
rect 169 337 170 338
rect 177 337 178 338
rect 178 337 179 338
rect 179 337 180 338
rect 180 337 181 338
rect 181 337 182 338
rect 182 337 183 338
rect 197 337 198 338
rect 198 337 199 338
rect 199 337 200 338
rect 288 337 289 338
rect 289 337 290 338
rect 300 337 301 338
rect 301 337 302 338
rect 302 337 303 338
rect 303 337 304 338
rect 340 337 341 338
rect 341 337 342 338
rect 342 337 343 338
rect 343 337 344 338
rect 344 337 345 338
rect 345 337 346 338
rect 346 337 347 338
rect 347 337 348 338
rect 348 337 349 338
rect 349 337 350 338
rect 350 337 351 338
rect 351 337 352 338
rect 352 337 353 338
rect 353 337 354 338
rect 354 337 355 338
rect 355 337 356 338
rect 356 337 357 338
rect 357 337 358 338
rect 358 337 359 338
rect 359 337 360 338
rect 360 337 361 338
rect 361 337 362 338
rect 362 337 363 338
rect 363 337 364 338
rect 364 337 365 338
rect 365 337 366 338
rect 366 337 367 338
rect 367 337 368 338
rect 368 337 369 338
rect 369 337 370 338
rect 370 337 371 338
rect 371 337 372 338
rect 372 337 373 338
rect 373 337 374 338
rect 374 337 375 338
rect 466 337 467 338
rect 467 337 468 338
rect 468 337 469 338
rect 469 337 470 338
rect 470 337 471 338
rect 471 337 472 338
rect 472 337 473 338
rect 473 337 474 338
rect 474 337 475 338
rect 475 337 476 338
rect 50 336 51 337
rect 51 336 52 337
rect 52 336 53 337
rect 53 336 54 337
rect 54 336 55 337
rect 55 336 56 337
rect 56 336 57 337
rect 57 336 58 337
rect 160 336 161 337
rect 161 336 162 337
rect 168 336 169 337
rect 169 336 170 337
rect 176 336 177 337
rect 177 336 178 337
rect 178 336 179 337
rect 179 336 180 337
rect 180 336 181 337
rect 181 336 182 337
rect 182 336 183 337
rect 287 336 288 337
rect 288 336 289 337
rect 289 336 290 337
rect 290 336 291 337
rect 299 336 300 337
rect 300 336 301 337
rect 301 336 302 337
rect 302 336 303 337
rect 303 336 304 337
rect 310 336 311 337
rect 339 336 340 337
rect 340 336 341 337
rect 341 336 342 337
rect 342 336 343 337
rect 343 336 344 337
rect 344 336 345 337
rect 345 336 346 337
rect 346 336 347 337
rect 347 336 348 337
rect 348 336 349 337
rect 349 336 350 337
rect 350 336 351 337
rect 351 336 352 337
rect 352 336 353 337
rect 353 336 354 337
rect 354 336 355 337
rect 355 336 356 337
rect 356 336 357 337
rect 357 336 358 337
rect 358 336 359 337
rect 359 336 360 337
rect 360 336 361 337
rect 361 336 362 337
rect 362 336 363 337
rect 363 336 364 337
rect 364 336 365 337
rect 365 336 366 337
rect 366 336 367 337
rect 367 336 368 337
rect 368 336 369 337
rect 369 336 370 337
rect 370 336 371 337
rect 371 336 372 337
rect 372 336 373 337
rect 373 336 374 337
rect 374 336 375 337
rect 375 336 376 337
rect 465 336 466 337
rect 466 336 467 337
rect 467 336 468 337
rect 468 336 469 337
rect 469 336 470 337
rect 470 336 471 337
rect 471 336 472 337
rect 472 336 473 337
rect 473 336 474 337
rect 474 336 475 337
rect 49 335 50 336
rect 50 335 51 336
rect 51 335 52 336
rect 52 335 53 336
rect 53 335 54 336
rect 54 335 55 336
rect 55 335 56 336
rect 56 335 57 336
rect 57 335 58 336
rect 160 335 161 336
rect 161 335 162 336
rect 162 335 163 336
rect 167 335 168 336
rect 168 335 169 336
rect 169 335 170 336
rect 176 335 177 336
rect 177 335 178 336
rect 178 335 179 336
rect 179 335 180 336
rect 180 335 181 336
rect 181 335 182 336
rect 182 335 183 336
rect 287 335 288 336
rect 288 335 289 336
rect 289 335 290 336
rect 290 335 291 336
rect 298 335 299 336
rect 299 335 300 336
rect 300 335 301 336
rect 301 335 302 336
rect 302 335 303 336
rect 303 335 304 336
rect 309 335 310 336
rect 310 335 311 336
rect 339 335 340 336
rect 340 335 341 336
rect 341 335 342 336
rect 342 335 343 336
rect 343 335 344 336
rect 344 335 345 336
rect 345 335 346 336
rect 346 335 347 336
rect 347 335 348 336
rect 348 335 349 336
rect 349 335 350 336
rect 350 335 351 336
rect 351 335 352 336
rect 352 335 353 336
rect 353 335 354 336
rect 354 335 355 336
rect 355 335 356 336
rect 356 335 357 336
rect 357 335 358 336
rect 358 335 359 336
rect 359 335 360 336
rect 360 335 361 336
rect 361 335 362 336
rect 362 335 363 336
rect 363 335 364 336
rect 364 335 365 336
rect 365 335 366 336
rect 366 335 367 336
rect 367 335 368 336
rect 368 335 369 336
rect 369 335 370 336
rect 370 335 371 336
rect 371 335 372 336
rect 372 335 373 336
rect 373 335 374 336
rect 374 335 375 336
rect 375 335 376 336
rect 464 335 465 336
rect 465 335 466 336
rect 466 335 467 336
rect 467 335 468 336
rect 468 335 469 336
rect 469 335 470 336
rect 470 335 471 336
rect 471 335 472 336
rect 472 335 473 336
rect 473 335 474 336
rect 49 334 50 335
rect 50 334 51 335
rect 51 334 52 335
rect 52 334 53 335
rect 53 334 54 335
rect 54 334 55 335
rect 55 334 56 335
rect 56 334 57 335
rect 57 334 58 335
rect 160 334 161 335
rect 161 334 162 335
rect 162 334 163 335
rect 167 334 168 335
rect 168 334 169 335
rect 169 334 170 335
rect 174 334 175 335
rect 175 334 176 335
rect 176 334 177 335
rect 177 334 178 335
rect 178 334 179 335
rect 179 334 180 335
rect 180 334 181 335
rect 181 334 182 335
rect 182 334 183 335
rect 183 334 184 335
rect 286 334 287 335
rect 287 334 288 335
rect 288 334 289 335
rect 289 334 290 335
rect 290 334 291 335
rect 297 334 298 335
rect 298 334 299 335
rect 299 334 300 335
rect 300 334 301 335
rect 301 334 302 335
rect 302 334 303 335
rect 309 334 310 335
rect 310 334 311 335
rect 338 334 339 335
rect 339 334 340 335
rect 340 334 341 335
rect 341 334 342 335
rect 342 334 343 335
rect 343 334 344 335
rect 344 334 345 335
rect 345 334 346 335
rect 346 334 347 335
rect 347 334 348 335
rect 348 334 349 335
rect 349 334 350 335
rect 350 334 351 335
rect 351 334 352 335
rect 352 334 353 335
rect 353 334 354 335
rect 354 334 355 335
rect 355 334 356 335
rect 356 334 357 335
rect 357 334 358 335
rect 358 334 359 335
rect 359 334 360 335
rect 360 334 361 335
rect 361 334 362 335
rect 362 334 363 335
rect 363 334 364 335
rect 364 334 365 335
rect 365 334 366 335
rect 366 334 367 335
rect 367 334 368 335
rect 368 334 369 335
rect 369 334 370 335
rect 370 334 371 335
rect 371 334 372 335
rect 372 334 373 335
rect 373 334 374 335
rect 374 334 375 335
rect 375 334 376 335
rect 464 334 465 335
rect 465 334 466 335
rect 466 334 467 335
rect 467 334 468 335
rect 468 334 469 335
rect 469 334 470 335
rect 470 334 471 335
rect 471 334 472 335
rect 472 334 473 335
rect 473 334 474 335
rect 49 333 50 334
rect 50 333 51 334
rect 51 333 52 334
rect 52 333 53 334
rect 53 333 54 334
rect 54 333 55 334
rect 55 333 56 334
rect 56 333 57 334
rect 57 333 58 334
rect 160 333 161 334
rect 161 333 162 334
rect 162 333 163 334
rect 163 333 164 334
rect 167 333 168 334
rect 168 333 169 334
rect 169 333 170 334
rect 170 333 171 334
rect 173 333 174 334
rect 174 333 175 334
rect 175 333 176 334
rect 176 333 177 334
rect 177 333 178 334
rect 178 333 179 334
rect 179 333 180 334
rect 180 333 181 334
rect 181 333 182 334
rect 182 333 183 334
rect 183 333 184 334
rect 184 333 185 334
rect 285 333 286 334
rect 286 333 287 334
rect 287 333 288 334
rect 288 333 289 334
rect 289 333 290 334
rect 290 333 291 334
rect 297 333 298 334
rect 298 333 299 334
rect 299 333 300 334
rect 300 333 301 334
rect 301 333 302 334
rect 302 333 303 334
rect 307 333 308 334
rect 308 333 309 334
rect 309 333 310 334
rect 310 333 311 334
rect 338 333 339 334
rect 339 333 340 334
rect 340 333 341 334
rect 341 333 342 334
rect 342 333 343 334
rect 343 333 344 334
rect 344 333 345 334
rect 345 333 346 334
rect 346 333 347 334
rect 347 333 348 334
rect 348 333 349 334
rect 349 333 350 334
rect 350 333 351 334
rect 351 333 352 334
rect 352 333 353 334
rect 353 333 354 334
rect 354 333 355 334
rect 355 333 356 334
rect 356 333 357 334
rect 357 333 358 334
rect 358 333 359 334
rect 359 333 360 334
rect 360 333 361 334
rect 361 333 362 334
rect 362 333 363 334
rect 363 333 364 334
rect 364 333 365 334
rect 365 333 366 334
rect 366 333 367 334
rect 367 333 368 334
rect 368 333 369 334
rect 369 333 370 334
rect 370 333 371 334
rect 371 333 372 334
rect 372 333 373 334
rect 373 333 374 334
rect 374 333 375 334
rect 375 333 376 334
rect 463 333 464 334
rect 464 333 465 334
rect 465 333 466 334
rect 466 333 467 334
rect 467 333 468 334
rect 468 333 469 334
rect 469 333 470 334
rect 470 333 471 334
rect 471 333 472 334
rect 472 333 473 334
rect 49 332 50 333
rect 50 332 51 333
rect 51 332 52 333
rect 52 332 53 333
rect 53 332 54 333
rect 54 332 55 333
rect 55 332 56 333
rect 56 332 57 333
rect 57 332 58 333
rect 160 332 161 333
rect 161 332 162 333
rect 162 332 163 333
rect 163 332 164 333
rect 167 332 168 333
rect 168 332 169 333
rect 169 332 170 333
rect 170 332 171 333
rect 171 332 172 333
rect 172 332 173 333
rect 173 332 174 333
rect 174 332 175 333
rect 175 332 176 333
rect 176 332 177 333
rect 177 332 178 333
rect 178 332 179 333
rect 179 332 180 333
rect 180 332 181 333
rect 181 332 182 333
rect 182 332 183 333
rect 183 332 184 333
rect 184 332 185 333
rect 185 332 186 333
rect 285 332 286 333
rect 286 332 287 333
rect 287 332 288 333
rect 288 332 289 333
rect 289 332 290 333
rect 290 332 291 333
rect 296 332 297 333
rect 297 332 298 333
rect 298 332 299 333
rect 299 332 300 333
rect 300 332 301 333
rect 301 332 302 333
rect 302 332 303 333
rect 306 332 307 333
rect 307 332 308 333
rect 308 332 309 333
rect 309 332 310 333
rect 310 332 311 333
rect 337 332 338 333
rect 338 332 339 333
rect 339 332 340 333
rect 340 332 341 333
rect 341 332 342 333
rect 342 332 343 333
rect 343 332 344 333
rect 344 332 345 333
rect 345 332 346 333
rect 346 332 347 333
rect 347 332 348 333
rect 348 332 349 333
rect 349 332 350 333
rect 350 332 351 333
rect 351 332 352 333
rect 352 332 353 333
rect 353 332 354 333
rect 354 332 355 333
rect 355 332 356 333
rect 356 332 357 333
rect 357 332 358 333
rect 358 332 359 333
rect 359 332 360 333
rect 360 332 361 333
rect 361 332 362 333
rect 362 332 363 333
rect 363 332 364 333
rect 364 332 365 333
rect 365 332 366 333
rect 366 332 367 333
rect 367 332 368 333
rect 368 332 369 333
rect 369 332 370 333
rect 370 332 371 333
rect 371 332 372 333
rect 372 332 373 333
rect 373 332 374 333
rect 374 332 375 333
rect 375 332 376 333
rect 462 332 463 333
rect 463 332 464 333
rect 464 332 465 333
rect 465 332 466 333
rect 466 332 467 333
rect 467 332 468 333
rect 468 332 469 333
rect 469 332 470 333
rect 470 332 471 333
rect 471 332 472 333
rect 49 331 50 332
rect 50 331 51 332
rect 51 331 52 332
rect 52 331 53 332
rect 53 331 54 332
rect 54 331 55 332
rect 55 331 56 332
rect 56 331 57 332
rect 57 331 58 332
rect 149 331 150 332
rect 160 331 161 332
rect 161 331 162 332
rect 162 331 163 332
rect 163 331 164 332
rect 167 331 168 332
rect 168 331 169 332
rect 169 331 170 332
rect 170 331 171 332
rect 171 331 172 332
rect 172 331 173 332
rect 173 331 174 332
rect 174 331 175 332
rect 175 331 176 332
rect 176 331 177 332
rect 177 331 178 332
rect 178 331 179 332
rect 179 331 180 332
rect 180 331 181 332
rect 181 331 182 332
rect 182 331 183 332
rect 183 331 184 332
rect 184 331 185 332
rect 185 331 186 332
rect 284 331 285 332
rect 285 331 286 332
rect 286 331 287 332
rect 287 331 288 332
rect 288 331 289 332
rect 289 331 290 332
rect 290 331 291 332
rect 295 331 296 332
rect 296 331 297 332
rect 297 331 298 332
rect 298 331 299 332
rect 299 331 300 332
rect 300 331 301 332
rect 301 331 302 332
rect 305 331 306 332
rect 306 331 307 332
rect 307 331 308 332
rect 308 331 309 332
rect 309 331 310 332
rect 337 331 338 332
rect 338 331 339 332
rect 339 331 340 332
rect 340 331 341 332
rect 341 331 342 332
rect 342 331 343 332
rect 343 331 344 332
rect 344 331 345 332
rect 345 331 346 332
rect 346 331 347 332
rect 347 331 348 332
rect 348 331 349 332
rect 349 331 350 332
rect 350 331 351 332
rect 351 331 352 332
rect 352 331 353 332
rect 353 331 354 332
rect 354 331 355 332
rect 355 331 356 332
rect 356 331 357 332
rect 357 331 358 332
rect 358 331 359 332
rect 359 331 360 332
rect 360 331 361 332
rect 361 331 362 332
rect 362 331 363 332
rect 363 331 364 332
rect 364 331 365 332
rect 365 331 366 332
rect 366 331 367 332
rect 367 331 368 332
rect 368 331 369 332
rect 369 331 370 332
rect 370 331 371 332
rect 371 331 372 332
rect 372 331 373 332
rect 373 331 374 332
rect 374 331 375 332
rect 375 331 376 332
rect 461 331 462 332
rect 462 331 463 332
rect 463 331 464 332
rect 464 331 465 332
rect 465 331 466 332
rect 466 331 467 332
rect 467 331 468 332
rect 468 331 469 332
rect 469 331 470 332
rect 470 331 471 332
rect 49 330 50 331
rect 50 330 51 331
rect 51 330 52 331
rect 52 330 53 331
rect 53 330 54 331
rect 54 330 55 331
rect 55 330 56 331
rect 56 330 57 331
rect 149 330 150 331
rect 150 330 151 331
rect 161 330 162 331
rect 162 330 163 331
rect 163 330 164 331
rect 164 330 165 331
rect 167 330 168 331
rect 168 330 169 331
rect 169 330 170 331
rect 170 330 171 331
rect 171 330 172 331
rect 172 330 173 331
rect 173 330 174 331
rect 174 330 175 331
rect 175 330 176 331
rect 176 330 177 331
rect 182 330 183 331
rect 183 330 184 331
rect 184 330 185 331
rect 185 330 186 331
rect 186 330 187 331
rect 284 330 285 331
rect 285 330 286 331
rect 286 330 287 331
rect 287 330 288 331
rect 288 330 289 331
rect 289 330 290 331
rect 290 330 291 331
rect 294 330 295 331
rect 295 330 296 331
rect 296 330 297 331
rect 297 330 298 331
rect 298 330 299 331
rect 299 330 300 331
rect 300 330 301 331
rect 301 330 302 331
rect 303 330 304 331
rect 304 330 305 331
rect 305 330 306 331
rect 306 330 307 331
rect 307 330 308 331
rect 308 330 309 331
rect 309 330 310 331
rect 336 330 337 331
rect 337 330 338 331
rect 338 330 339 331
rect 339 330 340 331
rect 340 330 341 331
rect 341 330 342 331
rect 342 330 343 331
rect 343 330 344 331
rect 344 330 345 331
rect 345 330 346 331
rect 346 330 347 331
rect 347 330 348 331
rect 348 330 349 331
rect 349 330 350 331
rect 350 330 351 331
rect 351 330 352 331
rect 352 330 353 331
rect 353 330 354 331
rect 354 330 355 331
rect 355 330 356 331
rect 356 330 357 331
rect 357 330 358 331
rect 358 330 359 331
rect 359 330 360 331
rect 360 330 361 331
rect 361 330 362 331
rect 362 330 363 331
rect 363 330 364 331
rect 364 330 365 331
rect 365 330 366 331
rect 366 330 367 331
rect 367 330 368 331
rect 368 330 369 331
rect 369 330 370 331
rect 370 330 371 331
rect 371 330 372 331
rect 372 330 373 331
rect 373 330 374 331
rect 374 330 375 331
rect 375 330 376 331
rect 460 330 461 331
rect 461 330 462 331
rect 462 330 463 331
rect 463 330 464 331
rect 464 330 465 331
rect 465 330 466 331
rect 466 330 467 331
rect 467 330 468 331
rect 468 330 469 331
rect 469 330 470 331
rect 48 329 49 330
rect 49 329 50 330
rect 50 329 51 330
rect 51 329 52 330
rect 52 329 53 330
rect 53 329 54 330
rect 54 329 55 330
rect 55 329 56 330
rect 56 329 57 330
rect 150 329 151 330
rect 151 329 152 330
rect 161 329 162 330
rect 162 329 163 330
rect 163 329 164 330
rect 164 329 165 330
rect 167 329 168 330
rect 168 329 169 330
rect 169 329 170 330
rect 170 329 171 330
rect 171 329 172 330
rect 172 329 173 330
rect 173 329 174 330
rect 174 329 175 330
rect 184 329 185 330
rect 185 329 186 330
rect 186 329 187 330
rect 187 329 188 330
rect 283 329 284 330
rect 284 329 285 330
rect 285 329 286 330
rect 286 329 287 330
rect 287 329 288 330
rect 288 329 289 330
rect 289 329 290 330
rect 290 329 291 330
rect 293 329 294 330
rect 294 329 295 330
rect 295 329 296 330
rect 296 329 297 330
rect 297 329 298 330
rect 298 329 299 330
rect 299 329 300 330
rect 300 329 301 330
rect 301 329 302 330
rect 302 329 303 330
rect 303 329 304 330
rect 304 329 305 330
rect 305 329 306 330
rect 306 329 307 330
rect 307 329 308 330
rect 308 329 309 330
rect 309 329 310 330
rect 335 329 336 330
rect 336 329 337 330
rect 337 329 338 330
rect 338 329 339 330
rect 339 329 340 330
rect 340 329 341 330
rect 341 329 342 330
rect 342 329 343 330
rect 343 329 344 330
rect 344 329 345 330
rect 345 329 346 330
rect 346 329 347 330
rect 347 329 348 330
rect 348 329 349 330
rect 349 329 350 330
rect 350 329 351 330
rect 351 329 352 330
rect 352 329 353 330
rect 353 329 354 330
rect 354 329 355 330
rect 355 329 356 330
rect 356 329 357 330
rect 357 329 358 330
rect 358 329 359 330
rect 359 329 360 330
rect 360 329 361 330
rect 361 329 362 330
rect 362 329 363 330
rect 363 329 364 330
rect 364 329 365 330
rect 365 329 366 330
rect 366 329 367 330
rect 367 329 368 330
rect 368 329 369 330
rect 369 329 370 330
rect 370 329 371 330
rect 371 329 372 330
rect 372 329 373 330
rect 373 329 374 330
rect 374 329 375 330
rect 375 329 376 330
rect 459 329 460 330
rect 460 329 461 330
rect 461 329 462 330
rect 462 329 463 330
rect 463 329 464 330
rect 464 329 465 330
rect 465 329 466 330
rect 466 329 467 330
rect 467 329 468 330
rect 468 329 469 330
rect 48 328 49 329
rect 49 328 50 329
rect 50 328 51 329
rect 51 328 52 329
rect 52 328 53 329
rect 53 328 54 329
rect 54 328 55 329
rect 55 328 56 329
rect 56 328 57 329
rect 150 328 151 329
rect 151 328 152 329
rect 152 328 153 329
rect 161 328 162 329
rect 162 328 163 329
rect 163 328 164 329
rect 164 328 165 329
rect 165 328 166 329
rect 167 328 168 329
rect 168 328 169 329
rect 169 328 170 329
rect 170 328 171 329
rect 171 328 172 329
rect 172 328 173 329
rect 173 328 174 329
rect 174 328 175 329
rect 185 328 186 329
rect 186 328 187 329
rect 187 328 188 329
rect 188 328 189 329
rect 282 328 283 329
rect 283 328 284 329
rect 284 328 285 329
rect 285 328 286 329
rect 286 328 287 329
rect 287 328 288 329
rect 288 328 289 329
rect 289 328 290 329
rect 290 328 291 329
rect 291 328 292 329
rect 292 328 293 329
rect 293 328 294 329
rect 294 328 295 329
rect 295 328 296 329
rect 296 328 297 329
rect 297 328 298 329
rect 298 328 299 329
rect 299 328 300 329
rect 300 328 301 329
rect 301 328 302 329
rect 302 328 303 329
rect 303 328 304 329
rect 304 328 305 329
rect 305 328 306 329
rect 306 328 307 329
rect 307 328 308 329
rect 308 328 309 329
rect 334 328 335 329
rect 335 328 336 329
rect 336 328 337 329
rect 337 328 338 329
rect 338 328 339 329
rect 339 328 340 329
rect 340 328 341 329
rect 341 328 342 329
rect 342 328 343 329
rect 343 328 344 329
rect 344 328 345 329
rect 345 328 346 329
rect 346 328 347 329
rect 347 328 348 329
rect 348 328 349 329
rect 349 328 350 329
rect 350 328 351 329
rect 351 328 352 329
rect 352 328 353 329
rect 353 328 354 329
rect 354 328 355 329
rect 355 328 356 329
rect 356 328 357 329
rect 357 328 358 329
rect 358 328 359 329
rect 359 328 360 329
rect 360 328 361 329
rect 361 328 362 329
rect 362 328 363 329
rect 363 328 364 329
rect 364 328 365 329
rect 365 328 366 329
rect 366 328 367 329
rect 367 328 368 329
rect 368 328 369 329
rect 369 328 370 329
rect 370 328 371 329
rect 371 328 372 329
rect 372 328 373 329
rect 373 328 374 329
rect 374 328 375 329
rect 375 328 376 329
rect 458 328 459 329
rect 459 328 460 329
rect 460 328 461 329
rect 461 328 462 329
rect 462 328 463 329
rect 463 328 464 329
rect 464 328 465 329
rect 465 328 466 329
rect 466 328 467 329
rect 467 328 468 329
rect 48 327 49 328
rect 49 327 50 328
rect 50 327 51 328
rect 51 327 52 328
rect 52 327 53 328
rect 53 327 54 328
rect 54 327 55 328
rect 55 327 56 328
rect 56 327 57 328
rect 150 327 151 328
rect 151 327 152 328
rect 152 327 153 328
rect 153 327 154 328
rect 161 327 162 328
rect 162 327 163 328
rect 163 327 164 328
rect 164 327 165 328
rect 165 327 166 328
rect 166 327 167 328
rect 167 327 168 328
rect 168 327 169 328
rect 169 327 170 328
rect 170 327 171 328
rect 171 327 172 328
rect 172 327 173 328
rect 173 327 174 328
rect 187 327 188 328
rect 188 327 189 328
rect 282 327 283 328
rect 283 327 284 328
rect 284 327 285 328
rect 285 327 286 328
rect 286 327 287 328
rect 287 327 288 328
rect 288 327 289 328
rect 289 327 290 328
rect 290 327 291 328
rect 291 327 292 328
rect 292 327 293 328
rect 293 327 294 328
rect 294 327 295 328
rect 295 327 296 328
rect 296 327 297 328
rect 297 327 298 328
rect 298 327 299 328
rect 299 327 300 328
rect 300 327 301 328
rect 301 327 302 328
rect 302 327 303 328
rect 303 327 304 328
rect 304 327 305 328
rect 305 327 306 328
rect 306 327 307 328
rect 307 327 308 328
rect 334 327 335 328
rect 335 327 336 328
rect 336 327 337 328
rect 337 327 338 328
rect 338 327 339 328
rect 339 327 340 328
rect 340 327 341 328
rect 341 327 342 328
rect 342 327 343 328
rect 344 327 345 328
rect 345 327 346 328
rect 346 327 347 328
rect 347 327 348 328
rect 348 327 349 328
rect 349 327 350 328
rect 350 327 351 328
rect 351 327 352 328
rect 352 327 353 328
rect 353 327 354 328
rect 354 327 355 328
rect 355 327 356 328
rect 356 327 357 328
rect 357 327 358 328
rect 358 327 359 328
rect 359 327 360 328
rect 360 327 361 328
rect 361 327 362 328
rect 362 327 363 328
rect 363 327 364 328
rect 364 327 365 328
rect 365 327 366 328
rect 366 327 367 328
rect 367 327 368 328
rect 368 327 369 328
rect 369 327 370 328
rect 370 327 371 328
rect 371 327 372 328
rect 372 327 373 328
rect 373 327 374 328
rect 374 327 375 328
rect 375 327 376 328
rect 457 327 458 328
rect 458 327 459 328
rect 459 327 460 328
rect 460 327 461 328
rect 461 327 462 328
rect 462 327 463 328
rect 463 327 464 328
rect 464 327 465 328
rect 465 327 466 328
rect 466 327 467 328
rect 48 326 49 327
rect 49 326 50 327
rect 50 326 51 327
rect 51 326 52 327
rect 52 326 53 327
rect 53 326 54 327
rect 54 326 55 327
rect 55 326 56 327
rect 56 326 57 327
rect 151 326 152 327
rect 152 326 153 327
rect 153 326 154 327
rect 154 326 155 327
rect 155 326 156 327
rect 161 326 162 327
rect 162 326 163 327
rect 163 326 164 327
rect 164 326 165 327
rect 165 326 166 327
rect 166 326 167 327
rect 167 326 168 327
rect 168 326 169 327
rect 169 326 170 327
rect 170 326 171 327
rect 171 326 172 327
rect 172 326 173 327
rect 188 326 189 327
rect 189 326 190 327
rect 281 326 282 327
rect 282 326 283 327
rect 283 326 284 327
rect 284 326 285 327
rect 285 326 286 327
rect 286 326 287 327
rect 287 326 288 327
rect 288 326 289 327
rect 289 326 290 327
rect 290 326 291 327
rect 291 326 292 327
rect 292 326 293 327
rect 293 326 294 327
rect 294 326 295 327
rect 295 326 296 327
rect 296 326 297 327
rect 297 326 298 327
rect 298 326 299 327
rect 299 326 300 327
rect 300 326 301 327
rect 301 326 302 327
rect 302 326 303 327
rect 303 326 304 327
rect 304 326 305 327
rect 305 326 306 327
rect 306 326 307 327
rect 333 326 334 327
rect 334 326 335 327
rect 335 326 336 327
rect 336 326 337 327
rect 337 326 338 327
rect 338 326 339 327
rect 339 326 340 327
rect 340 326 341 327
rect 341 326 342 327
rect 342 326 343 327
rect 344 326 345 327
rect 345 326 346 327
rect 346 326 347 327
rect 347 326 348 327
rect 348 326 349 327
rect 349 326 350 327
rect 350 326 351 327
rect 351 326 352 327
rect 352 326 353 327
rect 353 326 354 327
rect 354 326 355 327
rect 355 326 356 327
rect 356 326 357 327
rect 357 326 358 327
rect 358 326 359 327
rect 359 326 360 327
rect 360 326 361 327
rect 361 326 362 327
rect 362 326 363 327
rect 363 326 364 327
rect 364 326 365 327
rect 365 326 366 327
rect 366 326 367 327
rect 367 326 368 327
rect 368 326 369 327
rect 369 326 370 327
rect 370 326 371 327
rect 371 326 372 327
rect 372 326 373 327
rect 373 326 374 327
rect 374 326 375 327
rect 375 326 376 327
rect 456 326 457 327
rect 457 326 458 327
rect 458 326 459 327
rect 459 326 460 327
rect 460 326 461 327
rect 461 326 462 327
rect 462 326 463 327
rect 463 326 464 327
rect 464 326 465 327
rect 465 326 466 327
rect 466 326 467 327
rect 48 325 49 326
rect 49 325 50 326
rect 50 325 51 326
rect 51 325 52 326
rect 52 325 53 326
rect 53 325 54 326
rect 54 325 55 326
rect 55 325 56 326
rect 56 325 57 326
rect 152 325 153 326
rect 153 325 154 326
rect 154 325 155 326
rect 155 325 156 326
rect 156 325 157 326
rect 157 325 158 326
rect 162 325 163 326
rect 163 325 164 326
rect 164 325 165 326
rect 165 325 166 326
rect 166 325 167 326
rect 167 325 168 326
rect 168 325 169 326
rect 169 325 170 326
rect 170 325 171 326
rect 171 325 172 326
rect 172 325 173 326
rect 189 325 190 326
rect 280 325 281 326
rect 281 325 282 326
rect 282 325 283 326
rect 283 325 284 326
rect 284 325 285 326
rect 285 325 286 326
rect 286 325 287 326
rect 287 325 288 326
rect 288 325 289 326
rect 289 325 290 326
rect 290 325 291 326
rect 291 325 292 326
rect 292 325 293 326
rect 293 325 294 326
rect 294 325 295 326
rect 295 325 296 326
rect 296 325 297 326
rect 297 325 298 326
rect 298 325 299 326
rect 299 325 300 326
rect 300 325 301 326
rect 301 325 302 326
rect 302 325 303 326
rect 303 325 304 326
rect 304 325 305 326
rect 305 325 306 326
rect 306 325 307 326
rect 332 325 333 326
rect 333 325 334 326
rect 334 325 335 326
rect 335 325 336 326
rect 336 325 337 326
rect 337 325 338 326
rect 338 325 339 326
rect 339 325 340 326
rect 340 325 341 326
rect 341 325 342 326
rect 344 325 345 326
rect 345 325 346 326
rect 346 325 347 326
rect 347 325 348 326
rect 348 325 349 326
rect 349 325 350 326
rect 350 325 351 326
rect 351 325 352 326
rect 352 325 353 326
rect 353 325 354 326
rect 354 325 355 326
rect 355 325 356 326
rect 356 325 357 326
rect 357 325 358 326
rect 358 325 359 326
rect 359 325 360 326
rect 360 325 361 326
rect 361 325 362 326
rect 362 325 363 326
rect 363 325 364 326
rect 364 325 365 326
rect 365 325 366 326
rect 366 325 367 326
rect 367 325 368 326
rect 368 325 369 326
rect 369 325 370 326
rect 370 325 371 326
rect 371 325 372 326
rect 372 325 373 326
rect 373 325 374 326
rect 374 325 375 326
rect 455 325 456 326
rect 456 325 457 326
rect 457 325 458 326
rect 458 325 459 326
rect 459 325 460 326
rect 460 325 461 326
rect 461 325 462 326
rect 462 325 463 326
rect 463 325 464 326
rect 464 325 465 326
rect 465 325 466 326
rect 48 324 49 325
rect 49 324 50 325
rect 50 324 51 325
rect 51 324 52 325
rect 52 324 53 325
rect 53 324 54 325
rect 54 324 55 325
rect 55 324 56 325
rect 56 324 57 325
rect 152 324 153 325
rect 153 324 154 325
rect 154 324 155 325
rect 155 324 156 325
rect 156 324 157 325
rect 157 324 158 325
rect 158 324 159 325
rect 159 324 160 325
rect 160 324 161 325
rect 161 324 162 325
rect 162 324 163 325
rect 163 324 164 325
rect 164 324 165 325
rect 165 324 166 325
rect 166 324 167 325
rect 167 324 168 325
rect 168 324 169 325
rect 169 324 170 325
rect 170 324 171 325
rect 171 324 172 325
rect 172 324 173 325
rect 279 324 280 325
rect 280 324 281 325
rect 281 324 282 325
rect 282 324 283 325
rect 283 324 284 325
rect 284 324 285 325
rect 285 324 286 325
rect 286 324 287 325
rect 287 324 288 325
rect 288 324 289 325
rect 289 324 290 325
rect 290 324 291 325
rect 291 324 292 325
rect 292 324 293 325
rect 293 324 294 325
rect 294 324 295 325
rect 295 324 296 325
rect 296 324 297 325
rect 297 324 298 325
rect 298 324 299 325
rect 299 324 300 325
rect 300 324 301 325
rect 301 324 302 325
rect 302 324 303 325
rect 303 324 304 325
rect 304 324 305 325
rect 331 324 332 325
rect 332 324 333 325
rect 333 324 334 325
rect 334 324 335 325
rect 335 324 336 325
rect 336 324 337 325
rect 337 324 338 325
rect 338 324 339 325
rect 339 324 340 325
rect 340 324 341 325
rect 344 324 345 325
rect 345 324 346 325
rect 346 324 347 325
rect 347 324 348 325
rect 348 324 349 325
rect 349 324 350 325
rect 350 324 351 325
rect 351 324 352 325
rect 352 324 353 325
rect 353 324 354 325
rect 354 324 355 325
rect 355 324 356 325
rect 356 324 357 325
rect 357 324 358 325
rect 358 324 359 325
rect 359 324 360 325
rect 360 324 361 325
rect 361 324 362 325
rect 362 324 363 325
rect 363 324 364 325
rect 364 324 365 325
rect 365 324 366 325
rect 366 324 367 325
rect 367 324 368 325
rect 368 324 369 325
rect 369 324 370 325
rect 370 324 371 325
rect 371 324 372 325
rect 372 324 373 325
rect 373 324 374 325
rect 374 324 375 325
rect 454 324 455 325
rect 455 324 456 325
rect 456 324 457 325
rect 457 324 458 325
rect 458 324 459 325
rect 459 324 460 325
rect 460 324 461 325
rect 461 324 462 325
rect 462 324 463 325
rect 463 324 464 325
rect 464 324 465 325
rect 48 323 49 324
rect 49 323 50 324
rect 50 323 51 324
rect 51 323 52 324
rect 52 323 53 324
rect 53 323 54 324
rect 54 323 55 324
rect 55 323 56 324
rect 153 323 154 324
rect 154 323 155 324
rect 155 323 156 324
rect 156 323 157 324
rect 157 323 158 324
rect 158 323 159 324
rect 159 323 160 324
rect 160 323 161 324
rect 161 323 162 324
rect 162 323 163 324
rect 163 323 164 324
rect 164 323 165 324
rect 165 323 166 324
rect 166 323 167 324
rect 167 323 168 324
rect 168 323 169 324
rect 169 323 170 324
rect 170 323 171 324
rect 171 323 172 324
rect 172 323 173 324
rect 279 323 280 324
rect 280 323 281 324
rect 281 323 282 324
rect 282 323 283 324
rect 283 323 284 324
rect 284 323 285 324
rect 285 323 286 324
rect 286 323 287 324
rect 287 323 288 324
rect 288 323 289 324
rect 289 323 290 324
rect 290 323 291 324
rect 291 323 292 324
rect 292 323 293 324
rect 293 323 294 324
rect 294 323 295 324
rect 295 323 296 324
rect 296 323 297 324
rect 297 323 298 324
rect 298 323 299 324
rect 299 323 300 324
rect 300 323 301 324
rect 301 323 302 324
rect 302 323 303 324
rect 303 323 304 324
rect 330 323 331 324
rect 331 323 332 324
rect 332 323 333 324
rect 333 323 334 324
rect 334 323 335 324
rect 335 323 336 324
rect 336 323 337 324
rect 337 323 338 324
rect 338 323 339 324
rect 343 323 344 324
rect 344 323 345 324
rect 345 323 346 324
rect 346 323 347 324
rect 347 323 348 324
rect 348 323 349 324
rect 349 323 350 324
rect 350 323 351 324
rect 351 323 352 324
rect 352 323 353 324
rect 353 323 354 324
rect 354 323 355 324
rect 355 323 356 324
rect 356 323 357 324
rect 357 323 358 324
rect 358 323 359 324
rect 359 323 360 324
rect 360 323 361 324
rect 361 323 362 324
rect 362 323 363 324
rect 363 323 364 324
rect 364 323 365 324
rect 365 323 366 324
rect 366 323 367 324
rect 367 323 368 324
rect 368 323 369 324
rect 369 323 370 324
rect 370 323 371 324
rect 371 323 372 324
rect 372 323 373 324
rect 373 323 374 324
rect 374 323 375 324
rect 452 323 453 324
rect 453 323 454 324
rect 454 323 455 324
rect 455 323 456 324
rect 456 323 457 324
rect 457 323 458 324
rect 458 323 459 324
rect 459 323 460 324
rect 460 323 461 324
rect 461 323 462 324
rect 462 323 463 324
rect 463 323 464 324
rect 48 322 49 323
rect 49 322 50 323
rect 50 322 51 323
rect 51 322 52 323
rect 52 322 53 323
rect 53 322 54 323
rect 54 322 55 323
rect 55 322 56 323
rect 154 322 155 323
rect 155 322 156 323
rect 156 322 157 323
rect 157 322 158 323
rect 158 322 159 323
rect 159 322 160 323
rect 160 322 161 323
rect 161 322 162 323
rect 162 322 163 323
rect 163 322 164 323
rect 164 322 165 323
rect 165 322 166 323
rect 166 322 167 323
rect 167 322 168 323
rect 168 322 169 323
rect 169 322 170 323
rect 170 322 171 323
rect 171 322 172 323
rect 172 322 173 323
rect 173 322 174 323
rect 180 322 181 323
rect 266 322 267 323
rect 278 322 279 323
rect 279 322 280 323
rect 280 322 281 323
rect 281 322 282 323
rect 282 322 283 323
rect 283 322 284 323
rect 284 322 285 323
rect 285 322 286 323
rect 286 322 287 323
rect 287 322 288 323
rect 288 322 289 323
rect 289 322 290 323
rect 290 322 291 323
rect 291 322 292 323
rect 292 322 293 323
rect 293 322 294 323
rect 294 322 295 323
rect 295 322 296 323
rect 296 322 297 323
rect 297 322 298 323
rect 298 322 299 323
rect 299 322 300 323
rect 300 322 301 323
rect 301 322 302 323
rect 302 322 303 323
rect 329 322 330 323
rect 330 322 331 323
rect 331 322 332 323
rect 332 322 333 323
rect 333 322 334 323
rect 334 322 335 323
rect 335 322 336 323
rect 336 322 337 323
rect 343 322 344 323
rect 344 322 345 323
rect 345 322 346 323
rect 346 322 347 323
rect 347 322 348 323
rect 348 322 349 323
rect 349 322 350 323
rect 350 322 351 323
rect 351 322 352 323
rect 352 322 353 323
rect 353 322 354 323
rect 354 322 355 323
rect 355 322 356 323
rect 356 322 357 323
rect 357 322 358 323
rect 358 322 359 323
rect 359 322 360 323
rect 360 322 361 323
rect 361 322 362 323
rect 362 322 363 323
rect 363 322 364 323
rect 364 322 365 323
rect 365 322 366 323
rect 366 322 367 323
rect 367 322 368 323
rect 368 322 369 323
rect 369 322 370 323
rect 370 322 371 323
rect 371 322 372 323
rect 372 322 373 323
rect 373 322 374 323
rect 374 322 375 323
rect 451 322 452 323
rect 452 322 453 323
rect 453 322 454 323
rect 454 322 455 323
rect 455 322 456 323
rect 456 322 457 323
rect 457 322 458 323
rect 458 322 459 323
rect 459 322 460 323
rect 460 322 461 323
rect 461 322 462 323
rect 48 321 49 322
rect 49 321 50 322
rect 50 321 51 322
rect 51 321 52 322
rect 52 321 53 322
rect 53 321 54 322
rect 54 321 55 322
rect 55 321 56 322
rect 155 321 156 322
rect 156 321 157 322
rect 157 321 158 322
rect 158 321 159 322
rect 159 321 160 322
rect 160 321 161 322
rect 161 321 162 322
rect 162 321 163 322
rect 163 321 164 322
rect 164 321 165 322
rect 165 321 166 322
rect 166 321 167 322
rect 167 321 168 322
rect 168 321 169 322
rect 169 321 170 322
rect 170 321 171 322
rect 171 321 172 322
rect 172 321 173 322
rect 173 321 174 322
rect 180 321 181 322
rect 265 321 266 322
rect 266 321 267 322
rect 277 321 278 322
rect 278 321 279 322
rect 279 321 280 322
rect 280 321 281 322
rect 281 321 282 322
rect 282 321 283 322
rect 283 321 284 322
rect 284 321 285 322
rect 285 321 286 322
rect 286 321 287 322
rect 287 321 288 322
rect 288 321 289 322
rect 289 321 290 322
rect 290 321 291 322
rect 291 321 292 322
rect 292 321 293 322
rect 293 321 294 322
rect 294 321 295 322
rect 295 321 296 322
rect 296 321 297 322
rect 297 321 298 322
rect 298 321 299 322
rect 299 321 300 322
rect 300 321 301 322
rect 301 321 302 322
rect 327 321 328 322
rect 328 321 329 322
rect 329 321 330 322
rect 330 321 331 322
rect 331 321 332 322
rect 332 321 333 322
rect 333 321 334 322
rect 342 321 343 322
rect 343 321 344 322
rect 344 321 345 322
rect 345 321 346 322
rect 346 321 347 322
rect 347 321 348 322
rect 348 321 349 322
rect 349 321 350 322
rect 350 321 351 322
rect 351 321 352 322
rect 352 321 353 322
rect 353 321 354 322
rect 354 321 355 322
rect 355 321 356 322
rect 356 321 357 322
rect 357 321 358 322
rect 358 321 359 322
rect 359 321 360 322
rect 360 321 361 322
rect 361 321 362 322
rect 362 321 363 322
rect 363 321 364 322
rect 364 321 365 322
rect 365 321 366 322
rect 366 321 367 322
rect 367 321 368 322
rect 368 321 369 322
rect 369 321 370 322
rect 370 321 371 322
rect 371 321 372 322
rect 372 321 373 322
rect 373 321 374 322
rect 374 321 375 322
rect 450 321 451 322
rect 451 321 452 322
rect 452 321 453 322
rect 453 321 454 322
rect 454 321 455 322
rect 455 321 456 322
rect 456 321 457 322
rect 457 321 458 322
rect 458 321 459 322
rect 459 321 460 322
rect 460 321 461 322
rect 48 320 49 321
rect 49 320 50 321
rect 50 320 51 321
rect 51 320 52 321
rect 52 320 53 321
rect 53 320 54 321
rect 54 320 55 321
rect 55 320 56 321
rect 156 320 157 321
rect 157 320 158 321
rect 158 320 159 321
rect 159 320 160 321
rect 160 320 161 321
rect 161 320 162 321
rect 162 320 163 321
rect 163 320 164 321
rect 164 320 165 321
rect 165 320 166 321
rect 166 320 167 321
rect 167 320 168 321
rect 168 320 169 321
rect 169 320 170 321
rect 170 320 171 321
rect 171 320 172 321
rect 172 320 173 321
rect 173 320 174 321
rect 174 320 175 321
rect 179 320 180 321
rect 180 320 181 321
rect 181 320 182 321
rect 264 320 265 321
rect 265 320 266 321
rect 266 320 267 321
rect 276 320 277 321
rect 277 320 278 321
rect 278 320 279 321
rect 279 320 280 321
rect 280 320 281 321
rect 281 320 282 321
rect 282 320 283 321
rect 283 320 284 321
rect 284 320 285 321
rect 285 320 286 321
rect 286 320 287 321
rect 287 320 288 321
rect 288 320 289 321
rect 289 320 290 321
rect 290 320 291 321
rect 291 320 292 321
rect 292 320 293 321
rect 293 320 294 321
rect 294 320 295 321
rect 295 320 296 321
rect 296 320 297 321
rect 297 320 298 321
rect 298 320 299 321
rect 299 320 300 321
rect 342 320 343 321
rect 343 320 344 321
rect 344 320 345 321
rect 345 320 346 321
rect 346 320 347 321
rect 347 320 348 321
rect 348 320 349 321
rect 349 320 350 321
rect 350 320 351 321
rect 351 320 352 321
rect 352 320 353 321
rect 353 320 354 321
rect 354 320 355 321
rect 355 320 356 321
rect 356 320 357 321
rect 357 320 358 321
rect 358 320 359 321
rect 359 320 360 321
rect 360 320 361 321
rect 361 320 362 321
rect 362 320 363 321
rect 363 320 364 321
rect 364 320 365 321
rect 365 320 366 321
rect 366 320 367 321
rect 367 320 368 321
rect 368 320 369 321
rect 369 320 370 321
rect 370 320 371 321
rect 371 320 372 321
rect 372 320 373 321
rect 373 320 374 321
rect 374 320 375 321
rect 449 320 450 321
rect 450 320 451 321
rect 451 320 452 321
rect 452 320 453 321
rect 453 320 454 321
rect 454 320 455 321
rect 455 320 456 321
rect 456 320 457 321
rect 457 320 458 321
rect 458 320 459 321
rect 459 320 460 321
rect 47 319 48 320
rect 48 319 49 320
rect 49 319 50 320
rect 50 319 51 320
rect 51 319 52 320
rect 52 319 53 320
rect 53 319 54 320
rect 54 319 55 320
rect 55 319 56 320
rect 157 319 158 320
rect 158 319 159 320
rect 159 319 160 320
rect 160 319 161 320
rect 161 319 162 320
rect 162 319 163 320
rect 163 319 164 320
rect 164 319 165 320
rect 165 319 166 320
rect 166 319 167 320
rect 167 319 168 320
rect 168 319 169 320
rect 169 319 170 320
rect 170 319 171 320
rect 171 319 172 320
rect 172 319 173 320
rect 173 319 174 320
rect 174 319 175 320
rect 175 319 176 320
rect 179 319 180 320
rect 180 319 181 320
rect 181 319 182 320
rect 263 319 264 320
rect 264 319 265 320
rect 265 319 266 320
rect 266 319 267 320
rect 275 319 276 320
rect 276 319 277 320
rect 277 319 278 320
rect 278 319 279 320
rect 279 319 280 320
rect 280 319 281 320
rect 281 319 282 320
rect 282 319 283 320
rect 283 319 284 320
rect 284 319 285 320
rect 285 319 286 320
rect 286 319 287 320
rect 287 319 288 320
rect 288 319 289 320
rect 289 319 290 320
rect 290 319 291 320
rect 291 319 292 320
rect 292 319 293 320
rect 293 319 294 320
rect 294 319 295 320
rect 295 319 296 320
rect 296 319 297 320
rect 297 319 298 320
rect 341 319 342 320
rect 342 319 343 320
rect 343 319 344 320
rect 344 319 345 320
rect 345 319 346 320
rect 346 319 347 320
rect 347 319 348 320
rect 348 319 349 320
rect 349 319 350 320
rect 350 319 351 320
rect 351 319 352 320
rect 352 319 353 320
rect 353 319 354 320
rect 354 319 355 320
rect 355 319 356 320
rect 356 319 357 320
rect 357 319 358 320
rect 358 319 359 320
rect 359 319 360 320
rect 360 319 361 320
rect 361 319 362 320
rect 362 319 363 320
rect 363 319 364 320
rect 364 319 365 320
rect 365 319 366 320
rect 366 319 367 320
rect 367 319 368 320
rect 368 319 369 320
rect 369 319 370 320
rect 370 319 371 320
rect 371 319 372 320
rect 372 319 373 320
rect 373 319 374 320
rect 448 319 449 320
rect 449 319 450 320
rect 450 319 451 320
rect 451 319 452 320
rect 452 319 453 320
rect 453 319 454 320
rect 454 319 455 320
rect 455 319 456 320
rect 456 319 457 320
rect 457 319 458 320
rect 458 319 459 320
rect 47 318 48 319
rect 48 318 49 319
rect 49 318 50 319
rect 50 318 51 319
rect 51 318 52 319
rect 52 318 53 319
rect 53 318 54 319
rect 54 318 55 319
rect 55 318 56 319
rect 159 318 160 319
rect 160 318 161 319
rect 161 318 162 319
rect 162 318 163 319
rect 163 318 164 319
rect 164 318 165 319
rect 165 318 166 319
rect 166 318 167 319
rect 167 318 168 319
rect 168 318 169 319
rect 169 318 170 319
rect 170 318 171 319
rect 171 318 172 319
rect 172 318 173 319
rect 173 318 174 319
rect 174 318 175 319
rect 175 318 176 319
rect 176 318 177 319
rect 179 318 180 319
rect 180 318 181 319
rect 181 318 182 319
rect 262 318 263 319
rect 263 318 264 319
rect 264 318 265 319
rect 265 318 266 319
rect 266 318 267 319
rect 273 318 274 319
rect 274 318 275 319
rect 275 318 276 319
rect 276 318 277 319
rect 277 318 278 319
rect 278 318 279 319
rect 279 318 280 319
rect 280 318 281 319
rect 281 318 282 319
rect 282 318 283 319
rect 283 318 284 319
rect 284 318 285 319
rect 285 318 286 319
rect 286 318 287 319
rect 287 318 288 319
rect 288 318 289 319
rect 289 318 290 319
rect 290 318 291 319
rect 291 318 292 319
rect 292 318 293 319
rect 293 318 294 319
rect 294 318 295 319
rect 295 318 296 319
rect 296 318 297 319
rect 341 318 342 319
rect 342 318 343 319
rect 343 318 344 319
rect 344 318 345 319
rect 345 318 346 319
rect 346 318 347 319
rect 347 318 348 319
rect 348 318 349 319
rect 349 318 350 319
rect 350 318 351 319
rect 351 318 352 319
rect 352 318 353 319
rect 353 318 354 319
rect 354 318 355 319
rect 355 318 356 319
rect 356 318 357 319
rect 357 318 358 319
rect 358 318 359 319
rect 359 318 360 319
rect 360 318 361 319
rect 361 318 362 319
rect 362 318 363 319
rect 363 318 364 319
rect 364 318 365 319
rect 365 318 366 319
rect 366 318 367 319
rect 367 318 368 319
rect 368 318 369 319
rect 369 318 370 319
rect 370 318 371 319
rect 371 318 372 319
rect 372 318 373 319
rect 373 318 374 319
rect 447 318 448 319
rect 448 318 449 319
rect 449 318 450 319
rect 450 318 451 319
rect 451 318 452 319
rect 452 318 453 319
rect 453 318 454 319
rect 454 318 455 319
rect 455 318 456 319
rect 456 318 457 319
rect 457 318 458 319
rect 47 317 48 318
rect 48 317 49 318
rect 49 317 50 318
rect 50 317 51 318
rect 51 317 52 318
rect 52 317 53 318
rect 53 317 54 318
rect 54 317 55 318
rect 55 317 56 318
rect 160 317 161 318
rect 161 317 162 318
rect 162 317 163 318
rect 163 317 164 318
rect 164 317 165 318
rect 165 317 166 318
rect 166 317 167 318
rect 167 317 168 318
rect 168 317 169 318
rect 169 317 170 318
rect 170 317 171 318
rect 171 317 172 318
rect 172 317 173 318
rect 173 317 174 318
rect 174 317 175 318
rect 175 317 176 318
rect 176 317 177 318
rect 177 317 178 318
rect 179 317 180 318
rect 180 317 181 318
rect 181 317 182 318
rect 182 317 183 318
rect 261 317 262 318
rect 262 317 263 318
rect 263 317 264 318
rect 264 317 265 318
rect 265 317 266 318
rect 266 317 267 318
rect 272 317 273 318
rect 273 317 274 318
rect 274 317 275 318
rect 275 317 276 318
rect 276 317 277 318
rect 277 317 278 318
rect 278 317 279 318
rect 279 317 280 318
rect 280 317 281 318
rect 281 317 282 318
rect 282 317 283 318
rect 283 317 284 318
rect 284 317 285 318
rect 285 317 286 318
rect 286 317 287 318
rect 287 317 288 318
rect 288 317 289 318
rect 289 317 290 318
rect 290 317 291 318
rect 291 317 292 318
rect 292 317 293 318
rect 293 317 294 318
rect 294 317 295 318
rect 340 317 341 318
rect 341 317 342 318
rect 342 317 343 318
rect 343 317 344 318
rect 344 317 345 318
rect 345 317 346 318
rect 346 317 347 318
rect 347 317 348 318
rect 348 317 349 318
rect 349 317 350 318
rect 350 317 351 318
rect 351 317 352 318
rect 352 317 353 318
rect 353 317 354 318
rect 354 317 355 318
rect 355 317 356 318
rect 356 317 357 318
rect 357 317 358 318
rect 358 317 359 318
rect 359 317 360 318
rect 360 317 361 318
rect 361 317 362 318
rect 362 317 363 318
rect 363 317 364 318
rect 364 317 365 318
rect 365 317 366 318
rect 366 317 367 318
rect 367 317 368 318
rect 368 317 369 318
rect 369 317 370 318
rect 370 317 371 318
rect 371 317 372 318
rect 372 317 373 318
rect 373 317 374 318
rect 445 317 446 318
rect 446 317 447 318
rect 447 317 448 318
rect 448 317 449 318
rect 449 317 450 318
rect 450 317 451 318
rect 451 317 452 318
rect 452 317 453 318
rect 453 317 454 318
rect 454 317 455 318
rect 455 317 456 318
rect 456 317 457 318
rect 47 316 48 317
rect 48 316 49 317
rect 49 316 50 317
rect 50 316 51 317
rect 51 316 52 317
rect 52 316 53 317
rect 53 316 54 317
rect 54 316 55 317
rect 55 316 56 317
rect 162 316 163 317
rect 163 316 164 317
rect 164 316 165 317
rect 165 316 166 317
rect 166 316 167 317
rect 167 316 168 317
rect 168 316 169 317
rect 169 316 170 317
rect 170 316 171 317
rect 171 316 172 317
rect 172 316 173 317
rect 173 316 174 317
rect 174 316 175 317
rect 175 316 176 317
rect 176 316 177 317
rect 177 316 178 317
rect 178 316 179 317
rect 179 316 180 317
rect 180 316 181 317
rect 181 316 182 317
rect 182 316 183 317
rect 261 316 262 317
rect 262 316 263 317
rect 263 316 264 317
rect 264 316 265 317
rect 265 316 266 317
rect 266 316 267 317
rect 267 316 268 317
rect 269 316 270 317
rect 270 316 271 317
rect 271 316 272 317
rect 272 316 273 317
rect 273 316 274 317
rect 274 316 275 317
rect 275 316 276 317
rect 276 316 277 317
rect 277 316 278 317
rect 278 316 279 317
rect 279 316 280 317
rect 280 316 281 317
rect 281 316 282 317
rect 282 316 283 317
rect 283 316 284 317
rect 284 316 285 317
rect 285 316 286 317
rect 286 316 287 317
rect 287 316 288 317
rect 288 316 289 317
rect 289 316 290 317
rect 290 316 291 317
rect 291 316 292 317
rect 340 316 341 317
rect 341 316 342 317
rect 342 316 343 317
rect 343 316 344 317
rect 344 316 345 317
rect 345 316 346 317
rect 346 316 347 317
rect 347 316 348 317
rect 348 316 349 317
rect 349 316 350 317
rect 350 316 351 317
rect 351 316 352 317
rect 352 316 353 317
rect 353 316 354 317
rect 354 316 355 317
rect 355 316 356 317
rect 356 316 357 317
rect 357 316 358 317
rect 358 316 359 317
rect 359 316 360 317
rect 360 316 361 317
rect 361 316 362 317
rect 362 316 363 317
rect 363 316 364 317
rect 364 316 365 317
rect 365 316 366 317
rect 366 316 367 317
rect 367 316 368 317
rect 368 316 369 317
rect 369 316 370 317
rect 370 316 371 317
rect 371 316 372 317
rect 372 316 373 317
rect 373 316 374 317
rect 444 316 445 317
rect 445 316 446 317
rect 446 316 447 317
rect 447 316 448 317
rect 448 316 449 317
rect 449 316 450 317
rect 450 316 451 317
rect 451 316 452 317
rect 452 316 453 317
rect 453 316 454 317
rect 454 316 455 317
rect 455 316 456 317
rect 47 315 48 316
rect 48 315 49 316
rect 49 315 50 316
rect 50 315 51 316
rect 51 315 52 316
rect 52 315 53 316
rect 53 315 54 316
rect 54 315 55 316
rect 55 315 56 316
rect 162 315 163 316
rect 163 315 164 316
rect 164 315 165 316
rect 165 315 166 316
rect 166 315 167 316
rect 167 315 168 316
rect 168 315 169 316
rect 169 315 170 316
rect 170 315 171 316
rect 171 315 172 316
rect 172 315 173 316
rect 173 315 174 316
rect 174 315 175 316
rect 175 315 176 316
rect 176 315 177 316
rect 177 315 178 316
rect 178 315 179 316
rect 179 315 180 316
rect 180 315 181 316
rect 181 315 182 316
rect 182 315 183 316
rect 260 315 261 316
rect 261 315 262 316
rect 262 315 263 316
rect 263 315 264 316
rect 264 315 265 316
rect 265 315 266 316
rect 266 315 267 316
rect 267 315 268 316
rect 268 315 269 316
rect 269 315 270 316
rect 270 315 271 316
rect 271 315 272 316
rect 272 315 273 316
rect 273 315 274 316
rect 274 315 275 316
rect 275 315 276 316
rect 276 315 277 316
rect 277 315 278 316
rect 278 315 279 316
rect 279 315 280 316
rect 280 315 281 316
rect 281 315 282 316
rect 282 315 283 316
rect 283 315 284 316
rect 284 315 285 316
rect 285 315 286 316
rect 286 315 287 316
rect 287 315 288 316
rect 288 315 289 316
rect 289 315 290 316
rect 339 315 340 316
rect 340 315 341 316
rect 341 315 342 316
rect 342 315 343 316
rect 343 315 344 316
rect 344 315 345 316
rect 345 315 346 316
rect 346 315 347 316
rect 347 315 348 316
rect 348 315 349 316
rect 349 315 350 316
rect 350 315 351 316
rect 351 315 352 316
rect 352 315 353 316
rect 353 315 354 316
rect 354 315 355 316
rect 355 315 356 316
rect 356 315 357 316
rect 357 315 358 316
rect 358 315 359 316
rect 359 315 360 316
rect 360 315 361 316
rect 361 315 362 316
rect 362 315 363 316
rect 363 315 364 316
rect 364 315 365 316
rect 365 315 366 316
rect 366 315 367 316
rect 367 315 368 316
rect 368 315 369 316
rect 369 315 370 316
rect 370 315 371 316
rect 371 315 372 316
rect 372 315 373 316
rect 443 315 444 316
rect 444 315 445 316
rect 445 315 446 316
rect 446 315 447 316
rect 447 315 448 316
rect 448 315 449 316
rect 449 315 450 316
rect 450 315 451 316
rect 451 315 452 316
rect 452 315 453 316
rect 453 315 454 316
rect 454 315 455 316
rect 47 314 48 315
rect 48 314 49 315
rect 49 314 50 315
rect 50 314 51 315
rect 51 314 52 315
rect 52 314 53 315
rect 53 314 54 315
rect 54 314 55 315
rect 55 314 56 315
rect 163 314 164 315
rect 164 314 165 315
rect 165 314 166 315
rect 166 314 167 315
rect 167 314 168 315
rect 168 314 169 315
rect 169 314 170 315
rect 170 314 171 315
rect 171 314 172 315
rect 172 314 173 315
rect 173 314 174 315
rect 174 314 175 315
rect 175 314 176 315
rect 176 314 177 315
rect 177 314 178 315
rect 178 314 179 315
rect 179 314 180 315
rect 180 314 181 315
rect 181 314 182 315
rect 182 314 183 315
rect 183 314 184 315
rect 259 314 260 315
rect 260 314 261 315
rect 261 314 262 315
rect 262 314 263 315
rect 263 314 264 315
rect 264 314 265 315
rect 265 314 266 315
rect 266 314 267 315
rect 267 314 268 315
rect 268 314 269 315
rect 269 314 270 315
rect 270 314 271 315
rect 271 314 272 315
rect 272 314 273 315
rect 273 314 274 315
rect 274 314 275 315
rect 275 314 276 315
rect 276 314 277 315
rect 277 314 278 315
rect 278 314 279 315
rect 279 314 280 315
rect 280 314 281 315
rect 281 314 282 315
rect 282 314 283 315
rect 283 314 284 315
rect 284 314 285 315
rect 285 314 286 315
rect 286 314 287 315
rect 287 314 288 315
rect 338 314 339 315
rect 339 314 340 315
rect 340 314 341 315
rect 341 314 342 315
rect 342 314 343 315
rect 343 314 344 315
rect 344 314 345 315
rect 345 314 346 315
rect 346 314 347 315
rect 347 314 348 315
rect 348 314 349 315
rect 349 314 350 315
rect 350 314 351 315
rect 351 314 352 315
rect 352 314 353 315
rect 353 314 354 315
rect 354 314 355 315
rect 355 314 356 315
rect 356 314 357 315
rect 357 314 358 315
rect 358 314 359 315
rect 359 314 360 315
rect 360 314 361 315
rect 361 314 362 315
rect 362 314 363 315
rect 363 314 364 315
rect 364 314 365 315
rect 365 314 366 315
rect 366 314 367 315
rect 367 314 368 315
rect 368 314 369 315
rect 369 314 370 315
rect 370 314 371 315
rect 371 314 372 315
rect 372 314 373 315
rect 441 314 442 315
rect 442 314 443 315
rect 443 314 444 315
rect 444 314 445 315
rect 445 314 446 315
rect 446 314 447 315
rect 447 314 448 315
rect 448 314 449 315
rect 449 314 450 315
rect 450 314 451 315
rect 451 314 452 315
rect 452 314 453 315
rect 453 314 454 315
rect 47 313 48 314
rect 48 313 49 314
rect 49 313 50 314
rect 50 313 51 314
rect 51 313 52 314
rect 52 313 53 314
rect 53 313 54 314
rect 54 313 55 314
rect 55 313 56 314
rect 163 313 164 314
rect 164 313 165 314
rect 165 313 166 314
rect 166 313 167 314
rect 167 313 168 314
rect 168 313 169 314
rect 169 313 170 314
rect 170 313 171 314
rect 171 313 172 314
rect 172 313 173 314
rect 173 313 174 314
rect 174 313 175 314
rect 175 313 176 314
rect 176 313 177 314
rect 177 313 178 314
rect 178 313 179 314
rect 179 313 180 314
rect 180 313 181 314
rect 181 313 182 314
rect 182 313 183 314
rect 183 313 184 314
rect 184 313 185 314
rect 259 313 260 314
rect 260 313 261 314
rect 261 313 262 314
rect 262 313 263 314
rect 263 313 264 314
rect 264 313 265 314
rect 265 313 266 314
rect 266 313 267 314
rect 267 313 268 314
rect 268 313 269 314
rect 269 313 270 314
rect 270 313 271 314
rect 271 313 272 314
rect 272 313 273 314
rect 273 313 274 314
rect 274 313 275 314
rect 275 313 276 314
rect 276 313 277 314
rect 277 313 278 314
rect 278 313 279 314
rect 279 313 280 314
rect 280 313 281 314
rect 281 313 282 314
rect 282 313 283 314
rect 283 313 284 314
rect 284 313 285 314
rect 285 313 286 314
rect 286 313 287 314
rect 338 313 339 314
rect 339 313 340 314
rect 340 313 341 314
rect 341 313 342 314
rect 342 313 343 314
rect 343 313 344 314
rect 344 313 345 314
rect 345 313 346 314
rect 346 313 347 314
rect 347 313 348 314
rect 348 313 349 314
rect 349 313 350 314
rect 350 313 351 314
rect 351 313 352 314
rect 352 313 353 314
rect 353 313 354 314
rect 354 313 355 314
rect 355 313 356 314
rect 356 313 357 314
rect 357 313 358 314
rect 358 313 359 314
rect 359 313 360 314
rect 360 313 361 314
rect 361 313 362 314
rect 362 313 363 314
rect 363 313 364 314
rect 364 313 365 314
rect 365 313 366 314
rect 366 313 367 314
rect 367 313 368 314
rect 368 313 369 314
rect 369 313 370 314
rect 370 313 371 314
rect 371 313 372 314
rect 372 313 373 314
rect 440 313 441 314
rect 441 313 442 314
rect 442 313 443 314
rect 443 313 444 314
rect 444 313 445 314
rect 445 313 446 314
rect 446 313 447 314
rect 447 313 448 314
rect 448 313 449 314
rect 449 313 450 314
rect 450 313 451 314
rect 451 313 452 314
rect 47 312 48 313
rect 48 312 49 313
rect 49 312 50 313
rect 50 312 51 313
rect 51 312 52 313
rect 52 312 53 313
rect 53 312 54 313
rect 54 312 55 313
rect 55 312 56 313
rect 163 312 164 313
rect 164 312 165 313
rect 165 312 166 313
rect 166 312 167 313
rect 167 312 168 313
rect 168 312 169 313
rect 169 312 170 313
rect 170 312 171 313
rect 171 312 172 313
rect 172 312 173 313
rect 173 312 174 313
rect 174 312 175 313
rect 175 312 176 313
rect 176 312 177 313
rect 177 312 178 313
rect 178 312 179 313
rect 179 312 180 313
rect 180 312 181 313
rect 181 312 182 313
rect 182 312 183 313
rect 183 312 184 313
rect 184 312 185 313
rect 258 312 259 313
rect 259 312 260 313
rect 260 312 261 313
rect 261 312 262 313
rect 262 312 263 313
rect 263 312 264 313
rect 264 312 265 313
rect 265 312 266 313
rect 266 312 267 313
rect 267 312 268 313
rect 268 312 269 313
rect 269 312 270 313
rect 270 312 271 313
rect 271 312 272 313
rect 272 312 273 313
rect 273 312 274 313
rect 274 312 275 313
rect 275 312 276 313
rect 276 312 277 313
rect 277 312 278 313
rect 278 312 279 313
rect 279 312 280 313
rect 280 312 281 313
rect 281 312 282 313
rect 282 312 283 313
rect 283 312 284 313
rect 284 312 285 313
rect 285 312 286 313
rect 337 312 338 313
rect 338 312 339 313
rect 339 312 340 313
rect 340 312 341 313
rect 341 312 342 313
rect 342 312 343 313
rect 343 312 344 313
rect 344 312 345 313
rect 345 312 346 313
rect 346 312 347 313
rect 347 312 348 313
rect 348 312 349 313
rect 349 312 350 313
rect 350 312 351 313
rect 351 312 352 313
rect 352 312 353 313
rect 353 312 354 313
rect 354 312 355 313
rect 355 312 356 313
rect 356 312 357 313
rect 357 312 358 313
rect 358 312 359 313
rect 359 312 360 313
rect 360 312 361 313
rect 361 312 362 313
rect 362 312 363 313
rect 363 312 364 313
rect 364 312 365 313
rect 365 312 366 313
rect 366 312 367 313
rect 367 312 368 313
rect 368 312 369 313
rect 369 312 370 313
rect 370 312 371 313
rect 371 312 372 313
rect 439 312 440 313
rect 440 312 441 313
rect 441 312 442 313
rect 442 312 443 313
rect 443 312 444 313
rect 444 312 445 313
rect 445 312 446 313
rect 446 312 447 313
rect 447 312 448 313
rect 448 312 449 313
rect 449 312 450 313
rect 450 312 451 313
rect 47 311 48 312
rect 48 311 49 312
rect 49 311 50 312
rect 50 311 51 312
rect 51 311 52 312
rect 52 311 53 312
rect 53 311 54 312
rect 54 311 55 312
rect 55 311 56 312
rect 163 311 164 312
rect 164 311 165 312
rect 165 311 166 312
rect 166 311 167 312
rect 167 311 168 312
rect 168 311 169 312
rect 169 311 170 312
rect 170 311 171 312
rect 172 311 173 312
rect 173 311 174 312
rect 174 311 175 312
rect 175 311 176 312
rect 176 311 177 312
rect 177 311 178 312
rect 178 311 179 312
rect 179 311 180 312
rect 180 311 181 312
rect 181 311 182 312
rect 182 311 183 312
rect 183 311 184 312
rect 184 311 185 312
rect 185 311 186 312
rect 257 311 258 312
rect 258 311 259 312
rect 259 311 260 312
rect 260 311 261 312
rect 261 311 262 312
rect 262 311 263 312
rect 263 311 264 312
rect 264 311 265 312
rect 265 311 266 312
rect 266 311 267 312
rect 267 311 268 312
rect 268 311 269 312
rect 269 311 270 312
rect 270 311 271 312
rect 271 311 272 312
rect 272 311 273 312
rect 273 311 274 312
rect 274 311 275 312
rect 275 311 276 312
rect 276 311 277 312
rect 277 311 278 312
rect 278 311 279 312
rect 279 311 280 312
rect 280 311 281 312
rect 281 311 282 312
rect 282 311 283 312
rect 283 311 284 312
rect 336 311 337 312
rect 337 311 338 312
rect 338 311 339 312
rect 339 311 340 312
rect 340 311 341 312
rect 341 311 342 312
rect 342 311 343 312
rect 343 311 344 312
rect 344 311 345 312
rect 345 311 346 312
rect 346 311 347 312
rect 347 311 348 312
rect 348 311 349 312
rect 349 311 350 312
rect 350 311 351 312
rect 351 311 352 312
rect 352 311 353 312
rect 353 311 354 312
rect 354 311 355 312
rect 355 311 356 312
rect 356 311 357 312
rect 357 311 358 312
rect 358 311 359 312
rect 359 311 360 312
rect 360 311 361 312
rect 361 311 362 312
rect 362 311 363 312
rect 363 311 364 312
rect 364 311 365 312
rect 365 311 366 312
rect 366 311 367 312
rect 367 311 368 312
rect 368 311 369 312
rect 369 311 370 312
rect 370 311 371 312
rect 371 311 372 312
rect 437 311 438 312
rect 438 311 439 312
rect 439 311 440 312
rect 440 311 441 312
rect 441 311 442 312
rect 442 311 443 312
rect 443 311 444 312
rect 444 311 445 312
rect 445 311 446 312
rect 446 311 447 312
rect 447 311 448 312
rect 448 311 449 312
rect 449 311 450 312
rect 47 310 48 311
rect 48 310 49 311
rect 49 310 50 311
rect 50 310 51 311
rect 51 310 52 311
rect 52 310 53 311
rect 53 310 54 311
rect 54 310 55 311
rect 55 310 56 311
rect 163 310 164 311
rect 164 310 165 311
rect 165 310 166 311
rect 166 310 167 311
rect 167 310 168 311
rect 168 310 169 311
rect 169 310 170 311
rect 170 310 171 311
rect 174 310 175 311
rect 175 310 176 311
rect 176 310 177 311
rect 177 310 178 311
rect 178 310 179 311
rect 179 310 180 311
rect 180 310 181 311
rect 181 310 182 311
rect 182 310 183 311
rect 183 310 184 311
rect 184 310 185 311
rect 185 310 186 311
rect 186 310 187 311
rect 222 310 223 311
rect 256 310 257 311
rect 257 310 258 311
rect 258 310 259 311
rect 259 310 260 311
rect 260 310 261 311
rect 261 310 262 311
rect 262 310 263 311
rect 263 310 264 311
rect 264 310 265 311
rect 265 310 266 311
rect 266 310 267 311
rect 267 310 268 311
rect 268 310 269 311
rect 269 310 270 311
rect 270 310 271 311
rect 271 310 272 311
rect 272 310 273 311
rect 273 310 274 311
rect 274 310 275 311
rect 275 310 276 311
rect 276 310 277 311
rect 277 310 278 311
rect 278 310 279 311
rect 279 310 280 311
rect 280 310 281 311
rect 281 310 282 311
rect 336 310 337 311
rect 337 310 338 311
rect 338 310 339 311
rect 339 310 340 311
rect 340 310 341 311
rect 341 310 342 311
rect 342 310 343 311
rect 343 310 344 311
rect 344 310 345 311
rect 345 310 346 311
rect 346 310 347 311
rect 347 310 348 311
rect 348 310 349 311
rect 349 310 350 311
rect 350 310 351 311
rect 351 310 352 311
rect 352 310 353 311
rect 353 310 354 311
rect 354 310 355 311
rect 355 310 356 311
rect 356 310 357 311
rect 357 310 358 311
rect 358 310 359 311
rect 359 310 360 311
rect 360 310 361 311
rect 361 310 362 311
rect 362 310 363 311
rect 363 310 364 311
rect 364 310 365 311
rect 365 310 366 311
rect 366 310 367 311
rect 367 310 368 311
rect 368 310 369 311
rect 369 310 370 311
rect 370 310 371 311
rect 371 310 372 311
rect 372 310 373 311
rect 373 310 374 311
rect 374 310 375 311
rect 375 310 376 311
rect 376 310 377 311
rect 436 310 437 311
rect 437 310 438 311
rect 438 310 439 311
rect 439 310 440 311
rect 440 310 441 311
rect 441 310 442 311
rect 442 310 443 311
rect 443 310 444 311
rect 444 310 445 311
rect 445 310 446 311
rect 446 310 447 311
rect 447 310 448 311
rect 448 310 449 311
rect 47 309 48 310
rect 48 309 49 310
rect 49 309 50 310
rect 50 309 51 310
rect 51 309 52 310
rect 52 309 53 310
rect 53 309 54 310
rect 54 309 55 310
rect 55 309 56 310
rect 163 309 164 310
rect 164 309 165 310
rect 165 309 166 310
rect 166 309 167 310
rect 167 309 168 310
rect 168 309 169 310
rect 169 309 170 310
rect 170 309 171 310
rect 176 309 177 310
rect 177 309 178 310
rect 178 309 179 310
rect 179 309 180 310
rect 180 309 181 310
rect 181 309 182 310
rect 182 309 183 310
rect 183 309 184 310
rect 184 309 185 310
rect 185 309 186 310
rect 186 309 187 310
rect 187 309 188 310
rect 220 309 221 310
rect 221 309 222 310
rect 222 309 223 310
rect 256 309 257 310
rect 257 309 258 310
rect 258 309 259 310
rect 259 309 260 310
rect 260 309 261 310
rect 261 309 262 310
rect 262 309 263 310
rect 263 309 264 310
rect 264 309 265 310
rect 265 309 266 310
rect 266 309 267 310
rect 267 309 268 310
rect 268 309 269 310
rect 269 309 270 310
rect 270 309 271 310
rect 271 309 272 310
rect 272 309 273 310
rect 273 309 274 310
rect 274 309 275 310
rect 275 309 276 310
rect 276 309 277 310
rect 277 309 278 310
rect 278 309 279 310
rect 279 309 280 310
rect 335 309 336 310
rect 336 309 337 310
rect 337 309 338 310
rect 338 309 339 310
rect 339 309 340 310
rect 340 309 341 310
rect 341 309 342 310
rect 342 309 343 310
rect 343 309 344 310
rect 344 309 345 310
rect 345 309 346 310
rect 346 309 347 310
rect 347 309 348 310
rect 348 309 349 310
rect 349 309 350 310
rect 350 309 351 310
rect 351 309 352 310
rect 352 309 353 310
rect 353 309 354 310
rect 354 309 355 310
rect 355 309 356 310
rect 356 309 357 310
rect 357 309 358 310
rect 358 309 359 310
rect 359 309 360 310
rect 360 309 361 310
rect 361 309 362 310
rect 362 309 363 310
rect 363 309 364 310
rect 364 309 365 310
rect 365 309 366 310
rect 366 309 367 310
rect 367 309 368 310
rect 368 309 369 310
rect 369 309 370 310
rect 370 309 371 310
rect 371 309 372 310
rect 372 309 373 310
rect 373 309 374 310
rect 374 309 375 310
rect 375 309 376 310
rect 376 309 377 310
rect 377 309 378 310
rect 378 309 379 310
rect 379 309 380 310
rect 380 309 381 310
rect 434 309 435 310
rect 435 309 436 310
rect 436 309 437 310
rect 437 309 438 310
rect 438 309 439 310
rect 439 309 440 310
rect 440 309 441 310
rect 441 309 442 310
rect 442 309 443 310
rect 443 309 444 310
rect 444 309 445 310
rect 445 309 446 310
rect 446 309 447 310
rect 47 308 48 309
rect 48 308 49 309
rect 49 308 50 309
rect 50 308 51 309
rect 51 308 52 309
rect 52 308 53 309
rect 53 308 54 309
rect 54 308 55 309
rect 55 308 56 309
rect 164 308 165 309
rect 165 308 166 309
rect 166 308 167 309
rect 167 308 168 309
rect 168 308 169 309
rect 169 308 170 309
rect 170 308 171 309
rect 171 308 172 309
rect 178 308 179 309
rect 179 308 180 309
rect 180 308 181 309
rect 181 308 182 309
rect 182 308 183 309
rect 183 308 184 309
rect 184 308 185 309
rect 185 308 186 309
rect 186 308 187 309
rect 187 308 188 309
rect 188 308 189 309
rect 219 308 220 309
rect 220 308 221 309
rect 221 308 222 309
rect 255 308 256 309
rect 256 308 257 309
rect 257 308 258 309
rect 258 308 259 309
rect 259 308 260 309
rect 260 308 261 309
rect 261 308 262 309
rect 262 308 263 309
rect 263 308 264 309
rect 264 308 265 309
rect 265 308 266 309
rect 266 308 267 309
rect 267 308 268 309
rect 268 308 269 309
rect 269 308 270 309
rect 270 308 271 309
rect 271 308 272 309
rect 272 308 273 309
rect 273 308 274 309
rect 274 308 275 309
rect 275 308 276 309
rect 334 308 335 309
rect 335 308 336 309
rect 336 308 337 309
rect 337 308 338 309
rect 338 308 339 309
rect 339 308 340 309
rect 340 308 341 309
rect 341 308 342 309
rect 342 308 343 309
rect 343 308 344 309
rect 344 308 345 309
rect 345 308 346 309
rect 346 308 347 309
rect 347 308 348 309
rect 348 308 349 309
rect 349 308 350 309
rect 350 308 351 309
rect 351 308 352 309
rect 352 308 353 309
rect 353 308 354 309
rect 354 308 355 309
rect 355 308 356 309
rect 356 308 357 309
rect 357 308 358 309
rect 358 308 359 309
rect 359 308 360 309
rect 360 308 361 309
rect 361 308 362 309
rect 362 308 363 309
rect 363 308 364 309
rect 364 308 365 309
rect 365 308 366 309
rect 366 308 367 309
rect 367 308 368 309
rect 368 308 369 309
rect 369 308 370 309
rect 370 308 371 309
rect 371 308 372 309
rect 372 308 373 309
rect 373 308 374 309
rect 374 308 375 309
rect 375 308 376 309
rect 376 308 377 309
rect 377 308 378 309
rect 378 308 379 309
rect 379 308 380 309
rect 380 308 381 309
rect 381 308 382 309
rect 382 308 383 309
rect 383 308 384 309
rect 433 308 434 309
rect 434 308 435 309
rect 435 308 436 309
rect 436 308 437 309
rect 437 308 438 309
rect 438 308 439 309
rect 439 308 440 309
rect 440 308 441 309
rect 441 308 442 309
rect 442 308 443 309
rect 443 308 444 309
rect 444 308 445 309
rect 445 308 446 309
rect 47 307 48 308
rect 48 307 49 308
rect 49 307 50 308
rect 50 307 51 308
rect 51 307 52 308
rect 52 307 53 308
rect 53 307 54 308
rect 54 307 55 308
rect 55 307 56 308
rect 164 307 165 308
rect 165 307 166 308
rect 166 307 167 308
rect 167 307 168 308
rect 168 307 169 308
rect 169 307 170 308
rect 170 307 171 308
rect 171 307 172 308
rect 179 307 180 308
rect 180 307 181 308
rect 181 307 182 308
rect 182 307 183 308
rect 183 307 184 308
rect 184 307 185 308
rect 185 307 186 308
rect 186 307 187 308
rect 187 307 188 308
rect 188 307 189 308
rect 189 307 190 308
rect 218 307 219 308
rect 219 307 220 308
rect 220 307 221 308
rect 221 307 222 308
rect 254 307 255 308
rect 255 307 256 308
rect 256 307 257 308
rect 257 307 258 308
rect 258 307 259 308
rect 259 307 260 308
rect 260 307 261 308
rect 261 307 262 308
rect 262 307 263 308
rect 263 307 264 308
rect 264 307 265 308
rect 265 307 266 308
rect 266 307 267 308
rect 267 307 268 308
rect 268 307 269 308
rect 269 307 270 308
rect 270 307 271 308
rect 271 307 272 308
rect 272 307 273 308
rect 333 307 334 308
rect 334 307 335 308
rect 335 307 336 308
rect 336 307 337 308
rect 337 307 338 308
rect 338 307 339 308
rect 339 307 340 308
rect 340 307 341 308
rect 341 307 342 308
rect 342 307 343 308
rect 343 307 344 308
rect 344 307 345 308
rect 345 307 346 308
rect 346 307 347 308
rect 347 307 348 308
rect 348 307 349 308
rect 349 307 350 308
rect 350 307 351 308
rect 351 307 352 308
rect 352 307 353 308
rect 353 307 354 308
rect 354 307 355 308
rect 355 307 356 308
rect 356 307 357 308
rect 357 307 358 308
rect 358 307 359 308
rect 359 307 360 308
rect 360 307 361 308
rect 361 307 362 308
rect 362 307 363 308
rect 363 307 364 308
rect 364 307 365 308
rect 365 307 366 308
rect 366 307 367 308
rect 367 307 368 308
rect 368 307 369 308
rect 369 307 370 308
rect 370 307 371 308
rect 371 307 372 308
rect 372 307 373 308
rect 373 307 374 308
rect 374 307 375 308
rect 375 307 376 308
rect 376 307 377 308
rect 377 307 378 308
rect 378 307 379 308
rect 379 307 380 308
rect 380 307 381 308
rect 381 307 382 308
rect 382 307 383 308
rect 383 307 384 308
rect 384 307 385 308
rect 385 307 386 308
rect 431 307 432 308
rect 432 307 433 308
rect 433 307 434 308
rect 434 307 435 308
rect 435 307 436 308
rect 436 307 437 308
rect 437 307 438 308
rect 438 307 439 308
rect 439 307 440 308
rect 440 307 441 308
rect 441 307 442 308
rect 442 307 443 308
rect 443 307 444 308
rect 444 307 445 308
rect 47 306 48 307
rect 48 306 49 307
rect 49 306 50 307
rect 50 306 51 307
rect 51 306 52 307
rect 52 306 53 307
rect 53 306 54 307
rect 54 306 55 307
rect 55 306 56 307
rect 164 306 165 307
rect 165 306 166 307
rect 166 306 167 307
rect 167 306 168 307
rect 168 306 169 307
rect 169 306 170 307
rect 170 306 171 307
rect 171 306 172 307
rect 172 306 173 307
rect 181 306 182 307
rect 182 306 183 307
rect 183 306 184 307
rect 184 306 185 307
rect 185 306 186 307
rect 186 306 187 307
rect 187 306 188 307
rect 188 306 189 307
rect 189 306 190 307
rect 190 306 191 307
rect 217 306 218 307
rect 218 306 219 307
rect 219 306 220 307
rect 220 306 221 307
rect 253 306 254 307
rect 254 306 255 307
rect 255 306 256 307
rect 256 306 257 307
rect 257 306 258 307
rect 258 306 259 307
rect 259 306 260 307
rect 260 306 261 307
rect 261 306 262 307
rect 262 306 263 307
rect 263 306 264 307
rect 264 306 265 307
rect 265 306 266 307
rect 266 306 267 307
rect 267 306 268 307
rect 268 306 269 307
rect 269 306 270 307
rect 270 306 271 307
rect 333 306 334 307
rect 334 306 335 307
rect 335 306 336 307
rect 336 306 337 307
rect 337 306 338 307
rect 338 306 339 307
rect 339 306 340 307
rect 340 306 341 307
rect 341 306 342 307
rect 342 306 343 307
rect 343 306 344 307
rect 344 306 345 307
rect 345 306 346 307
rect 346 306 347 307
rect 347 306 348 307
rect 348 306 349 307
rect 349 306 350 307
rect 350 306 351 307
rect 351 306 352 307
rect 352 306 353 307
rect 353 306 354 307
rect 354 306 355 307
rect 355 306 356 307
rect 356 306 357 307
rect 357 306 358 307
rect 358 306 359 307
rect 359 306 360 307
rect 360 306 361 307
rect 361 306 362 307
rect 362 306 363 307
rect 363 306 364 307
rect 364 306 365 307
rect 365 306 366 307
rect 366 306 367 307
rect 367 306 368 307
rect 368 306 369 307
rect 369 306 370 307
rect 370 306 371 307
rect 371 306 372 307
rect 372 306 373 307
rect 373 306 374 307
rect 374 306 375 307
rect 375 306 376 307
rect 376 306 377 307
rect 377 306 378 307
rect 378 306 379 307
rect 379 306 380 307
rect 380 306 381 307
rect 381 306 382 307
rect 382 306 383 307
rect 383 306 384 307
rect 384 306 385 307
rect 385 306 386 307
rect 386 306 387 307
rect 387 306 388 307
rect 430 306 431 307
rect 431 306 432 307
rect 432 306 433 307
rect 433 306 434 307
rect 434 306 435 307
rect 435 306 436 307
rect 436 306 437 307
rect 437 306 438 307
rect 438 306 439 307
rect 439 306 440 307
rect 440 306 441 307
rect 441 306 442 307
rect 442 306 443 307
rect 47 305 48 306
rect 48 305 49 306
rect 49 305 50 306
rect 50 305 51 306
rect 51 305 52 306
rect 52 305 53 306
rect 53 305 54 306
rect 54 305 55 306
rect 55 305 56 306
rect 165 305 166 306
rect 166 305 167 306
rect 167 305 168 306
rect 168 305 169 306
rect 169 305 170 306
rect 170 305 171 306
rect 171 305 172 306
rect 172 305 173 306
rect 182 305 183 306
rect 183 305 184 306
rect 184 305 185 306
rect 185 305 186 306
rect 186 305 187 306
rect 187 305 188 306
rect 188 305 189 306
rect 189 305 190 306
rect 190 305 191 306
rect 191 305 192 306
rect 192 305 193 306
rect 217 305 218 306
rect 218 305 219 306
rect 219 305 220 306
rect 220 305 221 306
rect 252 305 253 306
rect 253 305 254 306
rect 254 305 255 306
rect 255 305 256 306
rect 256 305 257 306
rect 257 305 258 306
rect 258 305 259 306
rect 259 305 260 306
rect 260 305 261 306
rect 261 305 262 306
rect 262 305 263 306
rect 263 305 264 306
rect 264 305 265 306
rect 265 305 266 306
rect 266 305 267 306
rect 267 305 268 306
rect 268 305 269 306
rect 332 305 333 306
rect 333 305 334 306
rect 334 305 335 306
rect 335 305 336 306
rect 336 305 337 306
rect 337 305 338 306
rect 338 305 339 306
rect 339 305 340 306
rect 340 305 341 306
rect 341 305 342 306
rect 342 305 343 306
rect 343 305 344 306
rect 344 305 345 306
rect 345 305 346 306
rect 346 305 347 306
rect 347 305 348 306
rect 348 305 349 306
rect 349 305 350 306
rect 350 305 351 306
rect 351 305 352 306
rect 352 305 353 306
rect 353 305 354 306
rect 354 305 355 306
rect 355 305 356 306
rect 356 305 357 306
rect 357 305 358 306
rect 358 305 359 306
rect 359 305 360 306
rect 360 305 361 306
rect 361 305 362 306
rect 362 305 363 306
rect 363 305 364 306
rect 364 305 365 306
rect 365 305 366 306
rect 366 305 367 306
rect 367 305 368 306
rect 368 305 369 306
rect 369 305 370 306
rect 370 305 371 306
rect 371 305 372 306
rect 372 305 373 306
rect 373 305 374 306
rect 374 305 375 306
rect 375 305 376 306
rect 376 305 377 306
rect 377 305 378 306
rect 378 305 379 306
rect 379 305 380 306
rect 380 305 381 306
rect 381 305 382 306
rect 382 305 383 306
rect 383 305 384 306
rect 384 305 385 306
rect 385 305 386 306
rect 386 305 387 306
rect 387 305 388 306
rect 388 305 389 306
rect 428 305 429 306
rect 429 305 430 306
rect 430 305 431 306
rect 431 305 432 306
rect 432 305 433 306
rect 433 305 434 306
rect 434 305 435 306
rect 435 305 436 306
rect 436 305 437 306
rect 437 305 438 306
rect 438 305 439 306
rect 439 305 440 306
rect 440 305 441 306
rect 441 305 442 306
rect 47 304 48 305
rect 48 304 49 305
rect 49 304 50 305
rect 50 304 51 305
rect 51 304 52 305
rect 52 304 53 305
rect 53 304 54 305
rect 54 304 55 305
rect 55 304 56 305
rect 165 304 166 305
rect 166 304 167 305
rect 167 304 168 305
rect 168 304 169 305
rect 169 304 170 305
rect 170 304 171 305
rect 171 304 172 305
rect 172 304 173 305
rect 173 304 174 305
rect 185 304 186 305
rect 186 304 187 305
rect 187 304 188 305
rect 188 304 189 305
rect 189 304 190 305
rect 190 304 191 305
rect 191 304 192 305
rect 192 304 193 305
rect 193 304 194 305
rect 217 304 218 305
rect 218 304 219 305
rect 219 304 220 305
rect 220 304 221 305
rect 250 304 251 305
rect 251 304 252 305
rect 252 304 253 305
rect 253 304 254 305
rect 254 304 255 305
rect 255 304 256 305
rect 256 304 257 305
rect 257 304 258 305
rect 258 304 259 305
rect 259 304 260 305
rect 260 304 261 305
rect 261 304 262 305
rect 262 304 263 305
rect 263 304 264 305
rect 264 304 265 305
rect 265 304 266 305
rect 266 304 267 305
rect 331 304 332 305
rect 332 304 333 305
rect 333 304 334 305
rect 334 304 335 305
rect 335 304 336 305
rect 337 304 338 305
rect 338 304 339 305
rect 339 304 340 305
rect 340 304 341 305
rect 341 304 342 305
rect 342 304 343 305
rect 343 304 344 305
rect 344 304 345 305
rect 345 304 346 305
rect 346 304 347 305
rect 347 304 348 305
rect 348 304 349 305
rect 349 304 350 305
rect 350 304 351 305
rect 351 304 352 305
rect 352 304 353 305
rect 353 304 354 305
rect 354 304 355 305
rect 355 304 356 305
rect 356 304 357 305
rect 357 304 358 305
rect 358 304 359 305
rect 359 304 360 305
rect 360 304 361 305
rect 361 304 362 305
rect 362 304 363 305
rect 363 304 364 305
rect 364 304 365 305
rect 365 304 366 305
rect 366 304 367 305
rect 367 304 368 305
rect 368 304 369 305
rect 369 304 370 305
rect 370 304 371 305
rect 371 304 372 305
rect 372 304 373 305
rect 373 304 374 305
rect 374 304 375 305
rect 375 304 376 305
rect 376 304 377 305
rect 377 304 378 305
rect 378 304 379 305
rect 379 304 380 305
rect 380 304 381 305
rect 381 304 382 305
rect 382 304 383 305
rect 383 304 384 305
rect 384 304 385 305
rect 385 304 386 305
rect 386 304 387 305
rect 387 304 388 305
rect 388 304 389 305
rect 389 304 390 305
rect 390 304 391 305
rect 427 304 428 305
rect 428 304 429 305
rect 429 304 430 305
rect 430 304 431 305
rect 431 304 432 305
rect 432 304 433 305
rect 433 304 434 305
rect 434 304 435 305
rect 435 304 436 305
rect 436 304 437 305
rect 437 304 438 305
rect 438 304 439 305
rect 439 304 440 305
rect 47 303 48 304
rect 48 303 49 304
rect 49 303 50 304
rect 50 303 51 304
rect 51 303 52 304
rect 52 303 53 304
rect 53 303 54 304
rect 54 303 55 304
rect 55 303 56 304
rect 166 303 167 304
rect 167 303 168 304
rect 168 303 169 304
rect 169 303 170 304
rect 170 303 171 304
rect 171 303 172 304
rect 172 303 173 304
rect 173 303 174 304
rect 174 303 175 304
rect 187 303 188 304
rect 188 303 189 304
rect 189 303 190 304
rect 190 303 191 304
rect 191 303 192 304
rect 192 303 193 304
rect 193 303 194 304
rect 194 303 195 304
rect 195 303 196 304
rect 216 303 217 304
rect 217 303 218 304
rect 218 303 219 304
rect 219 303 220 304
rect 247 303 248 304
rect 248 303 249 304
rect 249 303 250 304
rect 250 303 251 304
rect 251 303 252 304
rect 252 303 253 304
rect 253 303 254 304
rect 254 303 255 304
rect 255 303 256 304
rect 256 303 257 304
rect 257 303 258 304
rect 258 303 259 304
rect 259 303 260 304
rect 260 303 261 304
rect 261 303 262 304
rect 262 303 263 304
rect 263 303 264 304
rect 264 303 265 304
rect 296 303 297 304
rect 297 303 298 304
rect 298 303 299 304
rect 330 303 331 304
rect 331 303 332 304
rect 332 303 333 304
rect 333 303 334 304
rect 337 303 338 304
rect 338 303 339 304
rect 339 303 340 304
rect 340 303 341 304
rect 341 303 342 304
rect 342 303 343 304
rect 343 303 344 304
rect 344 303 345 304
rect 345 303 346 304
rect 346 303 347 304
rect 347 303 348 304
rect 348 303 349 304
rect 349 303 350 304
rect 350 303 351 304
rect 351 303 352 304
rect 352 303 353 304
rect 353 303 354 304
rect 354 303 355 304
rect 355 303 356 304
rect 356 303 357 304
rect 357 303 358 304
rect 358 303 359 304
rect 359 303 360 304
rect 360 303 361 304
rect 361 303 362 304
rect 362 303 363 304
rect 363 303 364 304
rect 364 303 365 304
rect 365 303 366 304
rect 366 303 367 304
rect 367 303 368 304
rect 368 303 369 304
rect 369 303 370 304
rect 380 303 381 304
rect 381 303 382 304
rect 382 303 383 304
rect 383 303 384 304
rect 384 303 385 304
rect 385 303 386 304
rect 386 303 387 304
rect 387 303 388 304
rect 388 303 389 304
rect 389 303 390 304
rect 390 303 391 304
rect 391 303 392 304
rect 425 303 426 304
rect 426 303 427 304
rect 427 303 428 304
rect 428 303 429 304
rect 429 303 430 304
rect 430 303 431 304
rect 431 303 432 304
rect 432 303 433 304
rect 433 303 434 304
rect 434 303 435 304
rect 435 303 436 304
rect 436 303 437 304
rect 437 303 438 304
rect 438 303 439 304
rect 47 302 48 303
rect 48 302 49 303
rect 49 302 50 303
rect 50 302 51 303
rect 51 302 52 303
rect 52 302 53 303
rect 53 302 54 303
rect 54 302 55 303
rect 55 302 56 303
rect 167 302 168 303
rect 168 302 169 303
rect 169 302 170 303
rect 170 302 171 303
rect 171 302 172 303
rect 172 302 173 303
rect 173 302 174 303
rect 174 302 175 303
rect 175 302 176 303
rect 191 302 192 303
rect 192 302 193 303
rect 193 302 194 303
rect 216 302 217 303
rect 217 302 218 303
rect 218 302 219 303
rect 219 302 220 303
rect 240 302 241 303
rect 241 302 242 303
rect 242 302 243 303
rect 243 302 244 303
rect 244 302 245 303
rect 245 302 246 303
rect 246 302 247 303
rect 247 302 248 303
rect 248 302 249 303
rect 249 302 250 303
rect 250 302 251 303
rect 251 302 252 303
rect 252 302 253 303
rect 253 302 254 303
rect 254 302 255 303
rect 255 302 256 303
rect 256 302 257 303
rect 257 302 258 303
rect 258 302 259 303
rect 259 302 260 303
rect 260 302 261 303
rect 261 302 262 303
rect 262 302 263 303
rect 263 302 264 303
rect 291 302 292 303
rect 292 302 293 303
rect 293 302 294 303
rect 294 302 295 303
rect 295 302 296 303
rect 296 302 297 303
rect 297 302 298 303
rect 298 302 299 303
rect 299 302 300 303
rect 300 302 301 303
rect 301 302 302 303
rect 330 302 331 303
rect 331 302 332 303
rect 337 302 338 303
rect 338 302 339 303
rect 339 302 340 303
rect 340 302 341 303
rect 341 302 342 303
rect 342 302 343 303
rect 343 302 344 303
rect 344 302 345 303
rect 345 302 346 303
rect 346 302 347 303
rect 347 302 348 303
rect 348 302 349 303
rect 349 302 350 303
rect 350 302 351 303
rect 351 302 352 303
rect 352 302 353 303
rect 353 302 354 303
rect 354 302 355 303
rect 355 302 356 303
rect 356 302 357 303
rect 357 302 358 303
rect 358 302 359 303
rect 359 302 360 303
rect 360 302 361 303
rect 361 302 362 303
rect 362 302 363 303
rect 363 302 364 303
rect 364 302 365 303
rect 365 302 366 303
rect 366 302 367 303
rect 383 302 384 303
rect 384 302 385 303
rect 385 302 386 303
rect 386 302 387 303
rect 387 302 388 303
rect 388 302 389 303
rect 389 302 390 303
rect 390 302 391 303
rect 391 302 392 303
rect 392 302 393 303
rect 423 302 424 303
rect 424 302 425 303
rect 425 302 426 303
rect 426 302 427 303
rect 427 302 428 303
rect 428 302 429 303
rect 429 302 430 303
rect 430 302 431 303
rect 431 302 432 303
rect 432 302 433 303
rect 433 302 434 303
rect 434 302 435 303
rect 435 302 436 303
rect 436 302 437 303
rect 47 301 48 302
rect 48 301 49 302
rect 49 301 50 302
rect 50 301 51 302
rect 51 301 52 302
rect 52 301 53 302
rect 53 301 54 302
rect 54 301 55 302
rect 55 301 56 302
rect 167 301 168 302
rect 168 301 169 302
rect 169 301 170 302
rect 170 301 171 302
rect 171 301 172 302
rect 172 301 173 302
rect 173 301 174 302
rect 174 301 175 302
rect 175 301 176 302
rect 176 301 177 302
rect 201 301 202 302
rect 202 301 203 302
rect 216 301 217 302
rect 217 301 218 302
rect 218 301 219 302
rect 219 301 220 302
rect 241 301 242 302
rect 242 301 243 302
rect 243 301 244 302
rect 244 301 245 302
rect 245 301 246 302
rect 246 301 247 302
rect 247 301 248 302
rect 248 301 249 302
rect 249 301 250 302
rect 250 301 251 302
rect 251 301 252 302
rect 252 301 253 302
rect 253 301 254 302
rect 254 301 255 302
rect 255 301 256 302
rect 256 301 257 302
rect 257 301 258 302
rect 258 301 259 302
rect 259 301 260 302
rect 260 301 261 302
rect 261 301 262 302
rect 262 301 263 302
rect 263 301 264 302
rect 287 301 288 302
rect 288 301 289 302
rect 289 301 290 302
rect 290 301 291 302
rect 291 301 292 302
rect 292 301 293 302
rect 293 301 294 302
rect 294 301 295 302
rect 295 301 296 302
rect 296 301 297 302
rect 297 301 298 302
rect 298 301 299 302
rect 299 301 300 302
rect 300 301 301 302
rect 301 301 302 302
rect 302 301 303 302
rect 337 301 338 302
rect 338 301 339 302
rect 339 301 340 302
rect 340 301 341 302
rect 341 301 342 302
rect 342 301 343 302
rect 343 301 344 302
rect 344 301 345 302
rect 345 301 346 302
rect 346 301 347 302
rect 347 301 348 302
rect 348 301 349 302
rect 349 301 350 302
rect 350 301 351 302
rect 351 301 352 302
rect 352 301 353 302
rect 353 301 354 302
rect 354 301 355 302
rect 355 301 356 302
rect 356 301 357 302
rect 357 301 358 302
rect 358 301 359 302
rect 359 301 360 302
rect 360 301 361 302
rect 361 301 362 302
rect 362 301 363 302
rect 363 301 364 302
rect 364 301 365 302
rect 384 301 385 302
rect 385 301 386 302
rect 386 301 387 302
rect 387 301 388 302
rect 388 301 389 302
rect 389 301 390 302
rect 390 301 391 302
rect 391 301 392 302
rect 392 301 393 302
rect 393 301 394 302
rect 422 301 423 302
rect 423 301 424 302
rect 424 301 425 302
rect 425 301 426 302
rect 426 301 427 302
rect 427 301 428 302
rect 428 301 429 302
rect 429 301 430 302
rect 430 301 431 302
rect 431 301 432 302
rect 432 301 433 302
rect 433 301 434 302
rect 434 301 435 302
rect 435 301 436 302
rect 48 300 49 301
rect 49 300 50 301
rect 50 300 51 301
rect 51 300 52 301
rect 52 300 53 301
rect 53 300 54 301
rect 54 300 55 301
rect 55 300 56 301
rect 168 300 169 301
rect 169 300 170 301
rect 170 300 171 301
rect 171 300 172 301
rect 172 300 173 301
rect 173 300 174 301
rect 174 300 175 301
rect 175 300 176 301
rect 176 300 177 301
rect 177 300 178 301
rect 201 300 202 301
rect 202 300 203 301
rect 203 300 204 301
rect 216 300 217 301
rect 217 300 218 301
rect 218 300 219 301
rect 219 300 220 301
rect 241 300 242 301
rect 242 300 243 301
rect 243 300 244 301
rect 244 300 245 301
rect 245 300 246 301
rect 246 300 247 301
rect 247 300 248 301
rect 248 300 249 301
rect 249 300 250 301
rect 250 300 251 301
rect 251 300 252 301
rect 252 300 253 301
rect 253 300 254 301
rect 254 300 255 301
rect 255 300 256 301
rect 256 300 257 301
rect 257 300 258 301
rect 258 300 259 301
rect 259 300 260 301
rect 260 300 261 301
rect 261 300 262 301
rect 262 300 263 301
rect 263 300 264 301
rect 264 300 265 301
rect 284 300 285 301
rect 285 300 286 301
rect 286 300 287 301
rect 287 300 288 301
rect 288 300 289 301
rect 289 300 290 301
rect 290 300 291 301
rect 291 300 292 301
rect 292 300 293 301
rect 293 300 294 301
rect 294 300 295 301
rect 295 300 296 301
rect 296 300 297 301
rect 297 300 298 301
rect 298 300 299 301
rect 299 300 300 301
rect 300 300 301 301
rect 301 300 302 301
rect 302 300 303 301
rect 303 300 304 301
rect 337 300 338 301
rect 338 300 339 301
rect 339 300 340 301
rect 340 300 341 301
rect 341 300 342 301
rect 342 300 343 301
rect 343 300 344 301
rect 344 300 345 301
rect 345 300 346 301
rect 346 300 347 301
rect 347 300 348 301
rect 348 300 349 301
rect 349 300 350 301
rect 350 300 351 301
rect 351 300 352 301
rect 352 300 353 301
rect 353 300 354 301
rect 354 300 355 301
rect 355 300 356 301
rect 356 300 357 301
rect 357 300 358 301
rect 358 300 359 301
rect 359 300 360 301
rect 360 300 361 301
rect 361 300 362 301
rect 362 300 363 301
rect 385 300 386 301
rect 386 300 387 301
rect 387 300 388 301
rect 388 300 389 301
rect 389 300 390 301
rect 390 300 391 301
rect 391 300 392 301
rect 392 300 393 301
rect 393 300 394 301
rect 420 300 421 301
rect 421 300 422 301
rect 422 300 423 301
rect 423 300 424 301
rect 424 300 425 301
rect 425 300 426 301
rect 426 300 427 301
rect 427 300 428 301
rect 428 300 429 301
rect 429 300 430 301
rect 430 300 431 301
rect 431 300 432 301
rect 432 300 433 301
rect 433 300 434 301
rect 48 299 49 300
rect 49 299 50 300
rect 50 299 51 300
rect 51 299 52 300
rect 52 299 53 300
rect 53 299 54 300
rect 54 299 55 300
rect 55 299 56 300
rect 168 299 169 300
rect 169 299 170 300
rect 170 299 171 300
rect 171 299 172 300
rect 172 299 173 300
rect 173 299 174 300
rect 174 299 175 300
rect 175 299 176 300
rect 176 299 177 300
rect 177 299 178 300
rect 178 299 179 300
rect 201 299 202 300
rect 202 299 203 300
rect 203 299 204 300
rect 215 299 216 300
rect 216 299 217 300
rect 217 299 218 300
rect 218 299 219 300
rect 219 299 220 300
rect 242 299 243 300
rect 243 299 244 300
rect 244 299 245 300
rect 245 299 246 300
rect 246 299 247 300
rect 247 299 248 300
rect 248 299 249 300
rect 249 299 250 300
rect 250 299 251 300
rect 251 299 252 300
rect 252 299 253 300
rect 253 299 254 300
rect 254 299 255 300
rect 255 299 256 300
rect 256 299 257 300
rect 257 299 258 300
rect 258 299 259 300
rect 259 299 260 300
rect 260 299 261 300
rect 261 299 262 300
rect 262 299 263 300
rect 263 299 264 300
rect 264 299 265 300
rect 265 299 266 300
rect 281 299 282 300
rect 282 299 283 300
rect 283 299 284 300
rect 284 299 285 300
rect 285 299 286 300
rect 286 299 287 300
rect 287 299 288 300
rect 288 299 289 300
rect 289 299 290 300
rect 290 299 291 300
rect 291 299 292 300
rect 292 299 293 300
rect 293 299 294 300
rect 294 299 295 300
rect 295 299 296 300
rect 296 299 297 300
rect 297 299 298 300
rect 298 299 299 300
rect 299 299 300 300
rect 300 299 301 300
rect 301 299 302 300
rect 302 299 303 300
rect 303 299 304 300
rect 304 299 305 300
rect 337 299 338 300
rect 338 299 339 300
rect 339 299 340 300
rect 340 299 341 300
rect 341 299 342 300
rect 342 299 343 300
rect 343 299 344 300
rect 344 299 345 300
rect 345 299 346 300
rect 346 299 347 300
rect 347 299 348 300
rect 348 299 349 300
rect 349 299 350 300
rect 350 299 351 300
rect 351 299 352 300
rect 352 299 353 300
rect 353 299 354 300
rect 354 299 355 300
rect 355 299 356 300
rect 356 299 357 300
rect 357 299 358 300
rect 358 299 359 300
rect 359 299 360 300
rect 360 299 361 300
rect 361 299 362 300
rect 386 299 387 300
rect 387 299 388 300
rect 388 299 389 300
rect 389 299 390 300
rect 390 299 391 300
rect 391 299 392 300
rect 392 299 393 300
rect 393 299 394 300
rect 394 299 395 300
rect 418 299 419 300
rect 419 299 420 300
rect 420 299 421 300
rect 421 299 422 300
rect 422 299 423 300
rect 423 299 424 300
rect 424 299 425 300
rect 425 299 426 300
rect 426 299 427 300
rect 427 299 428 300
rect 428 299 429 300
rect 429 299 430 300
rect 430 299 431 300
rect 431 299 432 300
rect 432 299 433 300
rect 48 298 49 299
rect 49 298 50 299
rect 50 298 51 299
rect 51 298 52 299
rect 52 298 53 299
rect 53 298 54 299
rect 54 298 55 299
rect 55 298 56 299
rect 169 298 170 299
rect 170 298 171 299
rect 171 298 172 299
rect 172 298 173 299
rect 173 298 174 299
rect 174 298 175 299
rect 175 298 176 299
rect 176 298 177 299
rect 177 298 178 299
rect 178 298 179 299
rect 179 298 180 299
rect 201 298 202 299
rect 202 298 203 299
rect 203 298 204 299
rect 204 298 205 299
rect 216 298 217 299
rect 217 298 218 299
rect 218 298 219 299
rect 219 298 220 299
rect 244 298 245 299
rect 245 298 246 299
rect 246 298 247 299
rect 247 298 248 299
rect 248 298 249 299
rect 249 298 250 299
rect 250 298 251 299
rect 251 298 252 299
rect 252 298 253 299
rect 253 298 254 299
rect 254 298 255 299
rect 255 298 256 299
rect 256 298 257 299
rect 257 298 258 299
rect 258 298 259 299
rect 259 298 260 299
rect 260 298 261 299
rect 261 298 262 299
rect 262 298 263 299
rect 263 298 264 299
rect 278 298 279 299
rect 279 298 280 299
rect 280 298 281 299
rect 281 298 282 299
rect 282 298 283 299
rect 283 298 284 299
rect 284 298 285 299
rect 285 298 286 299
rect 286 298 287 299
rect 287 298 288 299
rect 288 298 289 299
rect 289 298 290 299
rect 290 298 291 299
rect 291 298 292 299
rect 292 298 293 299
rect 293 298 294 299
rect 294 298 295 299
rect 295 298 296 299
rect 296 298 297 299
rect 297 298 298 299
rect 298 298 299 299
rect 299 298 300 299
rect 300 298 301 299
rect 301 298 302 299
rect 302 298 303 299
rect 303 298 304 299
rect 304 298 305 299
rect 337 298 338 299
rect 338 298 339 299
rect 339 298 340 299
rect 340 298 341 299
rect 341 298 342 299
rect 342 298 343 299
rect 343 298 344 299
rect 344 298 345 299
rect 345 298 346 299
rect 346 298 347 299
rect 347 298 348 299
rect 348 298 349 299
rect 349 298 350 299
rect 350 298 351 299
rect 351 298 352 299
rect 352 298 353 299
rect 353 298 354 299
rect 354 298 355 299
rect 355 298 356 299
rect 356 298 357 299
rect 357 298 358 299
rect 358 298 359 299
rect 359 298 360 299
rect 387 298 388 299
rect 388 298 389 299
rect 389 298 390 299
rect 390 298 391 299
rect 391 298 392 299
rect 392 298 393 299
rect 393 298 394 299
rect 394 298 395 299
rect 395 298 396 299
rect 416 298 417 299
rect 417 298 418 299
rect 418 298 419 299
rect 419 298 420 299
rect 420 298 421 299
rect 421 298 422 299
rect 422 298 423 299
rect 423 298 424 299
rect 424 298 425 299
rect 425 298 426 299
rect 426 298 427 299
rect 427 298 428 299
rect 428 298 429 299
rect 429 298 430 299
rect 430 298 431 299
rect 48 297 49 298
rect 49 297 50 298
rect 50 297 51 298
rect 51 297 52 298
rect 52 297 53 298
rect 53 297 54 298
rect 54 297 55 298
rect 55 297 56 298
rect 56 297 57 298
rect 170 297 171 298
rect 171 297 172 298
rect 172 297 173 298
rect 173 297 174 298
rect 174 297 175 298
rect 175 297 176 298
rect 176 297 177 298
rect 177 297 178 298
rect 178 297 179 298
rect 179 297 180 298
rect 180 297 181 298
rect 181 297 182 298
rect 202 297 203 298
rect 203 297 204 298
rect 204 297 205 298
rect 216 297 217 298
rect 217 297 218 298
rect 218 297 219 298
rect 219 297 220 298
rect 245 297 246 298
rect 246 297 247 298
rect 247 297 248 298
rect 248 297 249 298
rect 249 297 250 298
rect 250 297 251 298
rect 251 297 252 298
rect 252 297 253 298
rect 253 297 254 298
rect 254 297 255 298
rect 255 297 256 298
rect 256 297 257 298
rect 257 297 258 298
rect 258 297 259 298
rect 259 297 260 298
rect 260 297 261 298
rect 275 297 276 298
rect 276 297 277 298
rect 277 297 278 298
rect 278 297 279 298
rect 279 297 280 298
rect 280 297 281 298
rect 281 297 282 298
rect 282 297 283 298
rect 283 297 284 298
rect 284 297 285 298
rect 285 297 286 298
rect 286 297 287 298
rect 287 297 288 298
rect 288 297 289 298
rect 289 297 290 298
rect 290 297 291 298
rect 291 297 292 298
rect 292 297 293 298
rect 337 297 338 298
rect 338 297 339 298
rect 339 297 340 298
rect 340 297 341 298
rect 341 297 342 298
rect 342 297 343 298
rect 343 297 344 298
rect 344 297 345 298
rect 345 297 346 298
rect 346 297 347 298
rect 347 297 348 298
rect 348 297 349 298
rect 349 297 350 298
rect 350 297 351 298
rect 351 297 352 298
rect 352 297 353 298
rect 353 297 354 298
rect 354 297 355 298
rect 355 297 356 298
rect 356 297 357 298
rect 357 297 358 298
rect 358 297 359 298
rect 388 297 389 298
rect 389 297 390 298
rect 390 297 391 298
rect 391 297 392 298
rect 392 297 393 298
rect 393 297 394 298
rect 394 297 395 298
rect 395 297 396 298
rect 415 297 416 298
rect 416 297 417 298
rect 417 297 418 298
rect 418 297 419 298
rect 419 297 420 298
rect 420 297 421 298
rect 421 297 422 298
rect 422 297 423 298
rect 423 297 424 298
rect 424 297 425 298
rect 425 297 426 298
rect 426 297 427 298
rect 427 297 428 298
rect 428 297 429 298
rect 429 297 430 298
rect 48 296 49 297
rect 49 296 50 297
rect 50 296 51 297
rect 51 296 52 297
rect 52 296 53 297
rect 53 296 54 297
rect 54 296 55 297
rect 55 296 56 297
rect 56 296 57 297
rect 171 296 172 297
rect 172 296 173 297
rect 173 296 174 297
rect 174 296 175 297
rect 175 296 176 297
rect 176 296 177 297
rect 177 296 178 297
rect 178 296 179 297
rect 179 296 180 297
rect 180 296 181 297
rect 181 296 182 297
rect 182 296 183 297
rect 183 296 184 297
rect 202 296 203 297
rect 203 296 204 297
rect 204 296 205 297
rect 205 296 206 297
rect 216 296 217 297
rect 217 296 218 297
rect 218 296 219 297
rect 219 296 220 297
rect 248 296 249 297
rect 249 296 250 297
rect 250 296 251 297
rect 251 296 252 297
rect 252 296 253 297
rect 253 296 254 297
rect 254 296 255 297
rect 255 296 256 297
rect 256 296 257 297
rect 273 296 274 297
rect 274 296 275 297
rect 275 296 276 297
rect 276 296 277 297
rect 277 296 278 297
rect 278 296 279 297
rect 279 296 280 297
rect 280 296 281 297
rect 281 296 282 297
rect 282 296 283 297
rect 283 296 284 297
rect 284 296 285 297
rect 285 296 286 297
rect 286 296 287 297
rect 287 296 288 297
rect 288 296 289 297
rect 289 296 290 297
rect 337 296 338 297
rect 338 296 339 297
rect 339 296 340 297
rect 340 296 341 297
rect 341 296 342 297
rect 342 296 343 297
rect 343 296 344 297
rect 344 296 345 297
rect 345 296 346 297
rect 346 296 347 297
rect 347 296 348 297
rect 348 296 349 297
rect 349 296 350 297
rect 350 296 351 297
rect 351 296 352 297
rect 352 296 353 297
rect 353 296 354 297
rect 354 296 355 297
rect 355 296 356 297
rect 356 296 357 297
rect 357 296 358 297
rect 389 296 390 297
rect 390 296 391 297
rect 391 296 392 297
rect 392 296 393 297
rect 393 296 394 297
rect 394 296 395 297
rect 395 296 396 297
rect 396 296 397 297
rect 413 296 414 297
rect 414 296 415 297
rect 415 296 416 297
rect 416 296 417 297
rect 417 296 418 297
rect 418 296 419 297
rect 419 296 420 297
rect 420 296 421 297
rect 421 296 422 297
rect 422 296 423 297
rect 423 296 424 297
rect 424 296 425 297
rect 425 296 426 297
rect 426 296 427 297
rect 427 296 428 297
rect 48 295 49 296
rect 49 295 50 296
rect 50 295 51 296
rect 51 295 52 296
rect 52 295 53 296
rect 53 295 54 296
rect 54 295 55 296
rect 55 295 56 296
rect 56 295 57 296
rect 171 295 172 296
rect 172 295 173 296
rect 173 295 174 296
rect 174 295 175 296
rect 175 295 176 296
rect 176 295 177 296
rect 177 295 178 296
rect 178 295 179 296
rect 179 295 180 296
rect 180 295 181 296
rect 181 295 182 296
rect 182 295 183 296
rect 183 295 184 296
rect 184 295 185 296
rect 185 295 186 296
rect 186 295 187 296
rect 202 295 203 296
rect 203 295 204 296
rect 204 295 205 296
rect 205 295 206 296
rect 217 295 218 296
rect 218 295 219 296
rect 219 295 220 296
rect 271 295 272 296
rect 272 295 273 296
rect 273 295 274 296
rect 274 295 275 296
rect 275 295 276 296
rect 276 295 277 296
rect 277 295 278 296
rect 278 295 279 296
rect 279 295 280 296
rect 280 295 281 296
rect 281 295 282 296
rect 282 295 283 296
rect 283 295 284 296
rect 284 295 285 296
rect 285 295 286 296
rect 286 295 287 296
rect 287 295 288 296
rect 288 295 289 296
rect 289 295 290 296
rect 290 295 291 296
rect 337 295 338 296
rect 338 295 339 296
rect 339 295 340 296
rect 340 295 341 296
rect 341 295 342 296
rect 342 295 343 296
rect 343 295 344 296
rect 344 295 345 296
rect 345 295 346 296
rect 346 295 347 296
rect 347 295 348 296
rect 348 295 349 296
rect 349 295 350 296
rect 350 295 351 296
rect 351 295 352 296
rect 352 295 353 296
rect 353 295 354 296
rect 354 295 355 296
rect 355 295 356 296
rect 356 295 357 296
rect 389 295 390 296
rect 390 295 391 296
rect 391 295 392 296
rect 392 295 393 296
rect 393 295 394 296
rect 394 295 395 296
rect 395 295 396 296
rect 396 295 397 296
rect 411 295 412 296
rect 412 295 413 296
rect 413 295 414 296
rect 414 295 415 296
rect 415 295 416 296
rect 416 295 417 296
rect 417 295 418 296
rect 418 295 419 296
rect 419 295 420 296
rect 420 295 421 296
rect 421 295 422 296
rect 422 295 423 296
rect 423 295 424 296
rect 424 295 425 296
rect 425 295 426 296
rect 48 294 49 295
rect 49 294 50 295
rect 50 294 51 295
rect 51 294 52 295
rect 52 294 53 295
rect 53 294 54 295
rect 54 294 55 295
rect 55 294 56 295
rect 56 294 57 295
rect 172 294 173 295
rect 173 294 174 295
rect 174 294 175 295
rect 175 294 176 295
rect 176 294 177 295
rect 177 294 178 295
rect 178 294 179 295
rect 179 294 180 295
rect 180 294 181 295
rect 181 294 182 295
rect 182 294 183 295
rect 183 294 184 295
rect 184 294 185 295
rect 185 294 186 295
rect 186 294 187 295
rect 187 294 188 295
rect 188 294 189 295
rect 189 294 190 295
rect 190 294 191 295
rect 202 294 203 295
rect 203 294 204 295
rect 204 294 205 295
rect 205 294 206 295
rect 268 294 269 295
rect 269 294 270 295
rect 270 294 271 295
rect 271 294 272 295
rect 272 294 273 295
rect 273 294 274 295
rect 274 294 275 295
rect 275 294 276 295
rect 276 294 277 295
rect 277 294 278 295
rect 278 294 279 295
rect 279 294 280 295
rect 280 294 281 295
rect 281 294 282 295
rect 285 294 286 295
rect 286 294 287 295
rect 287 294 288 295
rect 288 294 289 295
rect 289 294 290 295
rect 290 294 291 295
rect 337 294 338 295
rect 338 294 339 295
rect 339 294 340 295
rect 340 294 341 295
rect 341 294 342 295
rect 342 294 343 295
rect 343 294 344 295
rect 344 294 345 295
rect 345 294 346 295
rect 346 294 347 295
rect 347 294 348 295
rect 348 294 349 295
rect 349 294 350 295
rect 350 294 351 295
rect 351 294 352 295
rect 352 294 353 295
rect 353 294 354 295
rect 354 294 355 295
rect 355 294 356 295
rect 356 294 357 295
rect 374 294 375 295
rect 375 294 376 295
rect 390 294 391 295
rect 391 294 392 295
rect 392 294 393 295
rect 393 294 394 295
rect 394 294 395 295
rect 395 294 396 295
rect 396 294 397 295
rect 397 294 398 295
rect 409 294 410 295
rect 410 294 411 295
rect 411 294 412 295
rect 412 294 413 295
rect 413 294 414 295
rect 414 294 415 295
rect 415 294 416 295
rect 416 294 417 295
rect 417 294 418 295
rect 418 294 419 295
rect 419 294 420 295
rect 420 294 421 295
rect 421 294 422 295
rect 422 294 423 295
rect 423 294 424 295
rect 424 294 425 295
rect 48 293 49 294
rect 49 293 50 294
rect 50 293 51 294
rect 51 293 52 294
rect 52 293 53 294
rect 53 293 54 294
rect 54 293 55 294
rect 55 293 56 294
rect 56 293 57 294
rect 173 293 174 294
rect 174 293 175 294
rect 175 293 176 294
rect 176 293 177 294
rect 177 293 178 294
rect 178 293 179 294
rect 179 293 180 294
rect 180 293 181 294
rect 181 293 182 294
rect 182 293 183 294
rect 183 293 184 294
rect 184 293 185 294
rect 185 293 186 294
rect 186 293 187 294
rect 187 293 188 294
rect 188 293 189 294
rect 189 293 190 294
rect 190 293 191 294
rect 191 293 192 294
rect 192 293 193 294
rect 193 293 194 294
rect 194 293 195 294
rect 195 293 196 294
rect 196 293 197 294
rect 197 293 198 294
rect 198 293 199 294
rect 199 293 200 294
rect 200 293 201 294
rect 201 293 202 294
rect 202 293 203 294
rect 203 293 204 294
rect 204 293 205 294
rect 205 293 206 294
rect 266 293 267 294
rect 267 293 268 294
rect 268 293 269 294
rect 269 293 270 294
rect 270 293 271 294
rect 271 293 272 294
rect 272 293 273 294
rect 273 293 274 294
rect 274 293 275 294
rect 275 293 276 294
rect 276 293 277 294
rect 277 293 278 294
rect 278 293 279 294
rect 279 293 280 294
rect 286 293 287 294
rect 287 293 288 294
rect 288 293 289 294
rect 289 293 290 294
rect 290 293 291 294
rect 291 293 292 294
rect 337 293 338 294
rect 338 293 339 294
rect 339 293 340 294
rect 340 293 341 294
rect 341 293 342 294
rect 342 293 343 294
rect 343 293 344 294
rect 344 293 345 294
rect 345 293 346 294
rect 346 293 347 294
rect 347 293 348 294
rect 348 293 349 294
rect 349 293 350 294
rect 350 293 351 294
rect 351 293 352 294
rect 352 293 353 294
rect 353 293 354 294
rect 354 293 355 294
rect 355 293 356 294
rect 372 293 373 294
rect 373 293 374 294
rect 374 293 375 294
rect 375 293 376 294
rect 376 293 377 294
rect 390 293 391 294
rect 391 293 392 294
rect 392 293 393 294
rect 393 293 394 294
rect 394 293 395 294
rect 395 293 396 294
rect 396 293 397 294
rect 397 293 398 294
rect 407 293 408 294
rect 408 293 409 294
rect 409 293 410 294
rect 410 293 411 294
rect 411 293 412 294
rect 412 293 413 294
rect 413 293 414 294
rect 414 293 415 294
rect 415 293 416 294
rect 416 293 417 294
rect 417 293 418 294
rect 418 293 419 294
rect 419 293 420 294
rect 420 293 421 294
rect 421 293 422 294
rect 422 293 423 294
rect 49 292 50 293
rect 50 292 51 293
rect 51 292 52 293
rect 52 292 53 293
rect 53 292 54 293
rect 54 292 55 293
rect 55 292 56 293
rect 56 292 57 293
rect 173 292 174 293
rect 174 292 175 293
rect 175 292 176 293
rect 176 292 177 293
rect 177 292 178 293
rect 178 292 179 293
rect 179 292 180 293
rect 180 292 181 293
rect 181 292 182 293
rect 182 292 183 293
rect 183 292 184 293
rect 184 292 185 293
rect 185 292 186 293
rect 186 292 187 293
rect 187 292 188 293
rect 188 292 189 293
rect 189 292 190 293
rect 190 292 191 293
rect 191 292 192 293
rect 192 292 193 293
rect 193 292 194 293
rect 194 292 195 293
rect 195 292 196 293
rect 196 292 197 293
rect 197 292 198 293
rect 198 292 199 293
rect 199 292 200 293
rect 200 292 201 293
rect 201 292 202 293
rect 202 292 203 293
rect 203 292 204 293
rect 204 292 205 293
rect 264 292 265 293
rect 265 292 266 293
rect 266 292 267 293
rect 267 292 268 293
rect 268 292 269 293
rect 269 292 270 293
rect 270 292 271 293
rect 271 292 272 293
rect 272 292 273 293
rect 273 292 274 293
rect 274 292 275 293
rect 275 292 276 293
rect 276 292 277 293
rect 277 292 278 293
rect 278 292 279 293
rect 279 292 280 293
rect 286 292 287 293
rect 287 292 288 293
rect 288 292 289 293
rect 289 292 290 293
rect 290 292 291 293
rect 291 292 292 293
rect 337 292 338 293
rect 338 292 339 293
rect 339 292 340 293
rect 340 292 341 293
rect 341 292 342 293
rect 342 292 343 293
rect 343 292 344 293
rect 344 292 345 293
rect 345 292 346 293
rect 346 292 347 293
rect 347 292 348 293
rect 348 292 349 293
rect 349 292 350 293
rect 350 292 351 293
rect 351 292 352 293
rect 352 292 353 293
rect 353 292 354 293
rect 354 292 355 293
rect 355 292 356 293
rect 370 292 371 293
rect 371 292 372 293
rect 372 292 373 293
rect 373 292 374 293
rect 374 292 375 293
rect 375 292 376 293
rect 376 292 377 293
rect 377 292 378 293
rect 391 292 392 293
rect 392 292 393 293
rect 393 292 394 293
rect 394 292 395 293
rect 395 292 396 293
rect 396 292 397 293
rect 397 292 398 293
rect 405 292 406 293
rect 406 292 407 293
rect 407 292 408 293
rect 408 292 409 293
rect 409 292 410 293
rect 410 292 411 293
rect 411 292 412 293
rect 412 292 413 293
rect 413 292 414 293
rect 414 292 415 293
rect 415 292 416 293
rect 416 292 417 293
rect 417 292 418 293
rect 418 292 419 293
rect 419 292 420 293
rect 420 292 421 293
rect 49 291 50 292
rect 50 291 51 292
rect 51 291 52 292
rect 52 291 53 292
rect 53 291 54 292
rect 54 291 55 292
rect 55 291 56 292
rect 56 291 57 292
rect 57 291 58 292
rect 172 291 173 292
rect 173 291 174 292
rect 174 291 175 292
rect 175 291 176 292
rect 176 291 177 292
rect 177 291 178 292
rect 182 291 183 292
rect 183 291 184 292
rect 184 291 185 292
rect 185 291 186 292
rect 186 291 187 292
rect 187 291 188 292
rect 188 291 189 292
rect 189 291 190 292
rect 190 291 191 292
rect 191 291 192 292
rect 192 291 193 292
rect 193 291 194 292
rect 194 291 195 292
rect 195 291 196 292
rect 196 291 197 292
rect 197 291 198 292
rect 198 291 199 292
rect 199 291 200 292
rect 200 291 201 292
rect 201 291 202 292
rect 202 291 203 292
rect 203 291 204 292
rect 204 291 205 292
rect 262 291 263 292
rect 263 291 264 292
rect 264 291 265 292
rect 265 291 266 292
rect 266 291 267 292
rect 267 291 268 292
rect 268 291 269 292
rect 269 291 270 292
rect 270 291 271 292
rect 271 291 272 292
rect 272 291 273 292
rect 273 291 274 292
rect 274 291 275 292
rect 275 291 276 292
rect 276 291 277 292
rect 277 291 278 292
rect 278 291 279 292
rect 279 291 280 292
rect 287 291 288 292
rect 288 291 289 292
rect 289 291 290 292
rect 290 291 291 292
rect 291 291 292 292
rect 337 291 338 292
rect 338 291 339 292
rect 339 291 340 292
rect 340 291 341 292
rect 341 291 342 292
rect 342 291 343 292
rect 343 291 344 292
rect 344 291 345 292
rect 345 291 346 292
rect 346 291 347 292
rect 347 291 348 292
rect 348 291 349 292
rect 349 291 350 292
rect 350 291 351 292
rect 351 291 352 292
rect 352 291 353 292
rect 353 291 354 292
rect 354 291 355 292
rect 369 291 370 292
rect 370 291 371 292
rect 371 291 372 292
rect 372 291 373 292
rect 373 291 374 292
rect 374 291 375 292
rect 375 291 376 292
rect 376 291 377 292
rect 377 291 378 292
rect 391 291 392 292
rect 392 291 393 292
rect 393 291 394 292
rect 394 291 395 292
rect 395 291 396 292
rect 396 291 397 292
rect 397 291 398 292
rect 398 291 399 292
rect 402 291 403 292
rect 403 291 404 292
rect 404 291 405 292
rect 405 291 406 292
rect 406 291 407 292
rect 407 291 408 292
rect 408 291 409 292
rect 409 291 410 292
rect 410 291 411 292
rect 411 291 412 292
rect 412 291 413 292
rect 413 291 414 292
rect 414 291 415 292
rect 415 291 416 292
rect 416 291 417 292
rect 417 291 418 292
rect 418 291 419 292
rect 49 290 50 291
rect 50 290 51 291
rect 51 290 52 291
rect 52 290 53 291
rect 53 290 54 291
rect 54 290 55 291
rect 55 290 56 291
rect 56 290 57 291
rect 57 290 58 291
rect 172 290 173 291
rect 173 290 174 291
rect 174 290 175 291
rect 175 290 176 291
rect 176 290 177 291
rect 185 290 186 291
rect 186 290 187 291
rect 187 290 188 291
rect 188 290 189 291
rect 189 290 190 291
rect 190 290 191 291
rect 191 290 192 291
rect 192 290 193 291
rect 193 290 194 291
rect 194 290 195 291
rect 195 290 196 291
rect 196 290 197 291
rect 197 290 198 291
rect 198 290 199 291
rect 199 290 200 291
rect 200 290 201 291
rect 201 290 202 291
rect 202 290 203 291
rect 203 290 204 291
rect 259 290 260 291
rect 260 290 261 291
rect 261 290 262 291
rect 262 290 263 291
rect 263 290 264 291
rect 264 290 265 291
rect 265 290 266 291
rect 266 290 267 291
rect 267 290 268 291
rect 268 290 269 291
rect 269 290 270 291
rect 270 290 271 291
rect 271 290 272 291
rect 272 290 273 291
rect 273 290 274 291
rect 274 290 275 291
rect 275 290 276 291
rect 276 290 277 291
rect 277 290 278 291
rect 278 290 279 291
rect 279 290 280 291
rect 280 290 281 291
rect 287 290 288 291
rect 288 290 289 291
rect 289 290 290 291
rect 290 290 291 291
rect 291 290 292 291
rect 292 290 293 291
rect 337 290 338 291
rect 338 290 339 291
rect 339 290 340 291
rect 340 290 341 291
rect 341 290 342 291
rect 342 290 343 291
rect 343 290 344 291
rect 344 290 345 291
rect 345 290 346 291
rect 346 290 347 291
rect 347 290 348 291
rect 348 290 349 291
rect 349 290 350 291
rect 350 290 351 291
rect 351 290 352 291
rect 352 290 353 291
rect 353 290 354 291
rect 354 290 355 291
rect 367 290 368 291
rect 368 290 369 291
rect 369 290 370 291
rect 370 290 371 291
rect 371 290 372 291
rect 372 290 373 291
rect 373 290 374 291
rect 374 290 375 291
rect 375 290 376 291
rect 376 290 377 291
rect 377 290 378 291
rect 378 290 379 291
rect 391 290 392 291
rect 392 290 393 291
rect 393 290 394 291
rect 394 290 395 291
rect 395 290 396 291
rect 396 290 397 291
rect 397 290 398 291
rect 398 290 399 291
rect 400 290 401 291
rect 401 290 402 291
rect 402 290 403 291
rect 403 290 404 291
rect 404 290 405 291
rect 405 290 406 291
rect 406 290 407 291
rect 407 290 408 291
rect 408 290 409 291
rect 409 290 410 291
rect 410 290 411 291
rect 411 290 412 291
rect 412 290 413 291
rect 413 290 414 291
rect 414 290 415 291
rect 415 290 416 291
rect 416 290 417 291
rect 417 290 418 291
rect 49 289 50 290
rect 50 289 51 290
rect 51 289 52 290
rect 52 289 53 290
rect 53 289 54 290
rect 54 289 55 290
rect 55 289 56 290
rect 56 289 57 290
rect 57 289 58 290
rect 172 289 173 290
rect 173 289 174 290
rect 174 289 175 290
rect 175 289 176 290
rect 176 289 177 290
rect 187 289 188 290
rect 188 289 189 290
rect 189 289 190 290
rect 190 289 191 290
rect 191 289 192 290
rect 192 289 193 290
rect 193 289 194 290
rect 194 289 195 290
rect 195 289 196 290
rect 196 289 197 290
rect 197 289 198 290
rect 198 289 199 290
rect 199 289 200 290
rect 200 289 201 290
rect 201 289 202 290
rect 202 289 203 290
rect 203 289 204 290
rect 257 289 258 290
rect 258 289 259 290
rect 259 289 260 290
rect 260 289 261 290
rect 261 289 262 290
rect 262 289 263 290
rect 263 289 264 290
rect 264 289 265 290
rect 265 289 266 290
rect 266 289 267 290
rect 267 289 268 290
rect 268 289 269 290
rect 269 289 270 290
rect 270 289 271 290
rect 271 289 272 290
rect 272 289 273 290
rect 273 289 274 290
rect 274 289 275 290
rect 275 289 276 290
rect 276 289 277 290
rect 277 289 278 290
rect 278 289 279 290
rect 279 289 280 290
rect 280 289 281 290
rect 287 289 288 290
rect 288 289 289 290
rect 289 289 290 290
rect 290 289 291 290
rect 291 289 292 290
rect 292 289 293 290
rect 337 289 338 290
rect 338 289 339 290
rect 339 289 340 290
rect 340 289 341 290
rect 341 289 342 290
rect 342 289 343 290
rect 343 289 344 290
rect 344 289 345 290
rect 345 289 346 290
rect 346 289 347 290
rect 347 289 348 290
rect 348 289 349 290
rect 349 289 350 290
rect 350 289 351 290
rect 351 289 352 290
rect 352 289 353 290
rect 353 289 354 290
rect 354 289 355 290
rect 366 289 367 290
rect 367 289 368 290
rect 368 289 369 290
rect 369 289 370 290
rect 370 289 371 290
rect 371 289 372 290
rect 372 289 373 290
rect 373 289 374 290
rect 374 289 375 290
rect 375 289 376 290
rect 376 289 377 290
rect 377 289 378 290
rect 378 289 379 290
rect 391 289 392 290
rect 392 289 393 290
rect 393 289 394 290
rect 394 289 395 290
rect 395 289 396 290
rect 396 289 397 290
rect 397 289 398 290
rect 398 289 399 290
rect 399 289 400 290
rect 400 289 401 290
rect 401 289 402 290
rect 402 289 403 290
rect 403 289 404 290
rect 404 289 405 290
rect 405 289 406 290
rect 406 289 407 290
rect 407 289 408 290
rect 408 289 409 290
rect 409 289 410 290
rect 410 289 411 290
rect 411 289 412 290
rect 412 289 413 290
rect 413 289 414 290
rect 414 289 415 290
rect 415 289 416 290
rect 49 288 50 289
rect 50 288 51 289
rect 51 288 52 289
rect 52 288 53 289
rect 53 288 54 289
rect 54 288 55 289
rect 55 288 56 289
rect 56 288 57 289
rect 57 288 58 289
rect 172 288 173 289
rect 173 288 174 289
rect 174 288 175 289
rect 175 288 176 289
rect 176 288 177 289
rect 189 288 190 289
rect 190 288 191 289
rect 191 288 192 289
rect 192 288 193 289
rect 193 288 194 289
rect 194 288 195 289
rect 195 288 196 289
rect 196 288 197 289
rect 197 288 198 289
rect 198 288 199 289
rect 199 288 200 289
rect 200 288 201 289
rect 201 288 202 289
rect 202 288 203 289
rect 255 288 256 289
rect 256 288 257 289
rect 257 288 258 289
rect 258 288 259 289
rect 259 288 260 289
rect 260 288 261 289
rect 261 288 262 289
rect 262 288 263 289
rect 263 288 264 289
rect 264 288 265 289
rect 265 288 266 289
rect 266 288 267 289
rect 267 288 268 289
rect 268 288 269 289
rect 269 288 270 289
rect 270 288 271 289
rect 271 288 272 289
rect 272 288 273 289
rect 273 288 274 289
rect 274 288 275 289
rect 275 288 276 289
rect 276 288 277 289
rect 277 288 278 289
rect 278 288 279 289
rect 279 288 280 289
rect 280 288 281 289
rect 287 288 288 289
rect 288 288 289 289
rect 289 288 290 289
rect 290 288 291 289
rect 291 288 292 289
rect 292 288 293 289
rect 337 288 338 289
rect 338 288 339 289
rect 339 288 340 289
rect 340 288 341 289
rect 341 288 342 289
rect 342 288 343 289
rect 343 288 344 289
rect 344 288 345 289
rect 345 288 346 289
rect 346 288 347 289
rect 347 288 348 289
rect 348 288 349 289
rect 349 288 350 289
rect 350 288 351 289
rect 351 288 352 289
rect 352 288 353 289
rect 353 288 354 289
rect 365 288 366 289
rect 366 288 367 289
rect 367 288 368 289
rect 368 288 369 289
rect 369 288 370 289
rect 370 288 371 289
rect 371 288 372 289
rect 372 288 373 289
rect 373 288 374 289
rect 374 288 375 289
rect 375 288 376 289
rect 376 288 377 289
rect 377 288 378 289
rect 378 288 379 289
rect 379 288 380 289
rect 392 288 393 289
rect 393 288 394 289
rect 394 288 395 289
rect 395 288 396 289
rect 396 288 397 289
rect 397 288 398 289
rect 398 288 399 289
rect 399 288 400 289
rect 400 288 401 289
rect 401 288 402 289
rect 402 288 403 289
rect 403 288 404 289
rect 404 288 405 289
rect 405 288 406 289
rect 406 288 407 289
rect 407 288 408 289
rect 408 288 409 289
rect 409 288 410 289
rect 410 288 411 289
rect 411 288 412 289
rect 412 288 413 289
rect 413 288 414 289
rect 49 287 50 288
rect 50 287 51 288
rect 51 287 52 288
rect 52 287 53 288
rect 53 287 54 288
rect 54 287 55 288
rect 55 287 56 288
rect 56 287 57 288
rect 57 287 58 288
rect 171 287 172 288
rect 172 287 173 288
rect 173 287 174 288
rect 174 287 175 288
rect 175 287 176 288
rect 176 287 177 288
rect 186 287 187 288
rect 187 287 188 288
rect 188 287 189 288
rect 189 287 190 288
rect 190 287 191 288
rect 191 287 192 288
rect 192 287 193 288
rect 193 287 194 288
rect 194 287 195 288
rect 195 287 196 288
rect 196 287 197 288
rect 197 287 198 288
rect 198 287 199 288
rect 199 287 200 288
rect 200 287 201 288
rect 201 287 202 288
rect 252 287 253 288
rect 253 287 254 288
rect 254 287 255 288
rect 255 287 256 288
rect 256 287 257 288
rect 257 287 258 288
rect 258 287 259 288
rect 259 287 260 288
rect 260 287 261 288
rect 261 287 262 288
rect 262 287 263 288
rect 263 287 264 288
rect 264 287 265 288
rect 265 287 266 288
rect 266 287 267 288
rect 267 287 268 288
rect 268 287 269 288
rect 269 287 270 288
rect 270 287 271 288
rect 271 287 272 288
rect 272 287 273 288
rect 273 287 274 288
rect 274 287 275 288
rect 275 287 276 288
rect 276 287 277 288
rect 277 287 278 288
rect 278 287 279 288
rect 279 287 280 288
rect 280 287 281 288
rect 281 287 282 288
rect 288 287 289 288
rect 289 287 290 288
rect 290 287 291 288
rect 291 287 292 288
rect 292 287 293 288
rect 337 287 338 288
rect 338 287 339 288
rect 339 287 340 288
rect 340 287 341 288
rect 341 287 342 288
rect 342 287 343 288
rect 343 287 344 288
rect 344 287 345 288
rect 345 287 346 288
rect 346 287 347 288
rect 347 287 348 288
rect 348 287 349 288
rect 349 287 350 288
rect 350 287 351 288
rect 351 287 352 288
rect 352 287 353 288
rect 353 287 354 288
rect 364 287 365 288
rect 365 287 366 288
rect 366 287 367 288
rect 367 287 368 288
rect 368 287 369 288
rect 369 287 370 288
rect 370 287 371 288
rect 371 287 372 288
rect 372 287 373 288
rect 373 287 374 288
rect 374 287 375 288
rect 375 287 376 288
rect 376 287 377 288
rect 377 287 378 288
rect 378 287 379 288
rect 379 287 380 288
rect 392 287 393 288
rect 393 287 394 288
rect 394 287 395 288
rect 395 287 396 288
rect 396 287 397 288
rect 397 287 398 288
rect 398 287 399 288
rect 399 287 400 288
rect 400 287 401 288
rect 401 287 402 288
rect 402 287 403 288
rect 403 287 404 288
rect 404 287 405 288
rect 405 287 406 288
rect 406 287 407 288
rect 407 287 408 288
rect 408 287 409 288
rect 409 287 410 288
rect 410 287 411 288
rect 411 287 412 288
rect 50 286 51 287
rect 51 286 52 287
rect 52 286 53 287
rect 53 286 54 287
rect 54 286 55 287
rect 55 286 56 287
rect 56 286 57 287
rect 57 286 58 287
rect 58 286 59 287
rect 168 286 169 287
rect 169 286 170 287
rect 170 286 171 287
rect 171 286 172 287
rect 172 286 173 287
rect 173 286 174 287
rect 174 286 175 287
rect 175 286 176 287
rect 176 286 177 287
rect 186 286 187 287
rect 187 286 188 287
rect 188 286 189 287
rect 189 286 190 287
rect 190 286 191 287
rect 191 286 192 287
rect 192 286 193 287
rect 193 286 194 287
rect 194 286 195 287
rect 195 286 196 287
rect 196 286 197 287
rect 197 286 198 287
rect 198 286 199 287
rect 199 286 200 287
rect 200 286 201 287
rect 249 286 250 287
rect 250 286 251 287
rect 251 286 252 287
rect 252 286 253 287
rect 253 286 254 287
rect 254 286 255 287
rect 255 286 256 287
rect 256 286 257 287
rect 257 286 258 287
rect 258 286 259 287
rect 259 286 260 287
rect 260 286 261 287
rect 261 286 262 287
rect 262 286 263 287
rect 263 286 264 287
rect 264 286 265 287
rect 265 286 266 287
rect 266 286 267 287
rect 267 286 268 287
rect 269 286 270 287
rect 270 286 271 287
rect 271 286 272 287
rect 272 286 273 287
rect 273 286 274 287
rect 274 286 275 287
rect 275 286 276 287
rect 276 286 277 287
rect 277 286 278 287
rect 278 286 279 287
rect 279 286 280 287
rect 280 286 281 287
rect 281 286 282 287
rect 288 286 289 287
rect 289 286 290 287
rect 290 286 291 287
rect 291 286 292 287
rect 292 286 293 287
rect 337 286 338 287
rect 338 286 339 287
rect 339 286 340 287
rect 340 286 341 287
rect 341 286 342 287
rect 342 286 343 287
rect 343 286 344 287
rect 344 286 345 287
rect 345 286 346 287
rect 346 286 347 287
rect 347 286 348 287
rect 348 286 349 287
rect 349 286 350 287
rect 350 286 351 287
rect 351 286 352 287
rect 352 286 353 287
rect 353 286 354 287
rect 363 286 364 287
rect 364 286 365 287
rect 365 286 366 287
rect 366 286 367 287
rect 367 286 368 287
rect 368 286 369 287
rect 376 286 377 287
rect 377 286 378 287
rect 378 286 379 287
rect 379 286 380 287
rect 380 286 381 287
rect 392 286 393 287
rect 393 286 394 287
rect 394 286 395 287
rect 395 286 396 287
rect 396 286 397 287
rect 397 286 398 287
rect 398 286 399 287
rect 399 286 400 287
rect 400 286 401 287
rect 401 286 402 287
rect 402 286 403 287
rect 403 286 404 287
rect 404 286 405 287
rect 405 286 406 287
rect 406 286 407 287
rect 407 286 408 287
rect 408 286 409 287
rect 409 286 410 287
rect 50 285 51 286
rect 51 285 52 286
rect 52 285 53 286
rect 53 285 54 286
rect 54 285 55 286
rect 55 285 56 286
rect 56 285 57 286
rect 57 285 58 286
rect 58 285 59 286
rect 166 285 167 286
rect 167 285 168 286
rect 168 285 169 286
rect 169 285 170 286
rect 170 285 171 286
rect 171 285 172 286
rect 172 285 173 286
rect 173 285 174 286
rect 174 285 175 286
rect 175 285 176 286
rect 176 285 177 286
rect 186 285 187 286
rect 187 285 188 286
rect 188 285 189 286
rect 189 285 190 286
rect 190 285 191 286
rect 191 285 192 286
rect 192 285 193 286
rect 193 285 194 286
rect 194 285 195 286
rect 195 285 196 286
rect 196 285 197 286
rect 197 285 198 286
rect 198 285 199 286
rect 199 285 200 286
rect 237 285 238 286
rect 238 285 239 286
rect 239 285 240 286
rect 240 285 241 286
rect 241 285 242 286
rect 242 285 243 286
rect 243 285 244 286
rect 244 285 245 286
rect 245 285 246 286
rect 246 285 247 286
rect 247 285 248 286
rect 248 285 249 286
rect 249 285 250 286
rect 250 285 251 286
rect 251 285 252 286
rect 252 285 253 286
rect 253 285 254 286
rect 254 285 255 286
rect 255 285 256 286
rect 256 285 257 286
rect 257 285 258 286
rect 258 285 259 286
rect 259 285 260 286
rect 260 285 261 286
rect 261 285 262 286
rect 262 285 263 286
rect 263 285 264 286
rect 264 285 265 286
rect 265 285 266 286
rect 266 285 267 286
rect 270 285 271 286
rect 271 285 272 286
rect 272 285 273 286
rect 273 285 274 286
rect 274 285 275 286
rect 276 285 277 286
rect 277 285 278 286
rect 278 285 279 286
rect 279 285 280 286
rect 280 285 281 286
rect 281 285 282 286
rect 288 285 289 286
rect 289 285 290 286
rect 290 285 291 286
rect 291 285 292 286
rect 292 285 293 286
rect 337 285 338 286
rect 338 285 339 286
rect 339 285 340 286
rect 340 285 341 286
rect 341 285 342 286
rect 342 285 343 286
rect 343 285 344 286
rect 344 285 345 286
rect 345 285 346 286
rect 346 285 347 286
rect 347 285 348 286
rect 348 285 349 286
rect 349 285 350 286
rect 350 285 351 286
rect 351 285 352 286
rect 352 285 353 286
rect 353 285 354 286
rect 362 285 363 286
rect 363 285 364 286
rect 364 285 365 286
rect 365 285 366 286
rect 366 285 367 286
rect 367 285 368 286
rect 377 285 378 286
rect 378 285 379 286
rect 379 285 380 286
rect 380 285 381 286
rect 392 285 393 286
rect 393 285 394 286
rect 394 285 395 286
rect 395 285 396 286
rect 396 285 397 286
rect 397 285 398 286
rect 398 285 399 286
rect 399 285 400 286
rect 400 285 401 286
rect 401 285 402 286
rect 402 285 403 286
rect 403 285 404 286
rect 404 285 405 286
rect 405 285 406 286
rect 406 285 407 286
rect 407 285 408 286
rect 50 284 51 285
rect 51 284 52 285
rect 52 284 53 285
rect 53 284 54 285
rect 54 284 55 285
rect 55 284 56 285
rect 56 284 57 285
rect 57 284 58 285
rect 58 284 59 285
rect 164 284 165 285
rect 165 284 166 285
rect 166 284 167 285
rect 167 284 168 285
rect 168 284 169 285
rect 169 284 170 285
rect 170 284 171 285
rect 171 284 172 285
rect 172 284 173 285
rect 173 284 174 285
rect 174 284 175 285
rect 175 284 176 285
rect 176 284 177 285
rect 177 284 178 285
rect 187 284 188 285
rect 188 284 189 285
rect 189 284 190 285
rect 190 284 191 285
rect 191 284 192 285
rect 192 284 193 285
rect 193 284 194 285
rect 194 284 195 285
rect 195 284 196 285
rect 196 284 197 285
rect 197 284 198 285
rect 198 284 199 285
rect 237 284 238 285
rect 238 284 239 285
rect 239 284 240 285
rect 240 284 241 285
rect 241 284 242 285
rect 242 284 243 285
rect 243 284 244 285
rect 244 284 245 285
rect 245 284 246 285
rect 246 284 247 285
rect 247 284 248 285
rect 248 284 249 285
rect 249 284 250 285
rect 250 284 251 285
rect 251 284 252 285
rect 252 284 253 285
rect 253 284 254 285
rect 254 284 255 285
rect 255 284 256 285
rect 256 284 257 285
rect 257 284 258 285
rect 258 284 259 285
rect 259 284 260 285
rect 260 284 261 285
rect 263 284 264 285
rect 264 284 265 285
rect 265 284 266 285
rect 266 284 267 285
rect 267 284 268 285
rect 276 284 277 285
rect 277 284 278 285
rect 278 284 279 285
rect 279 284 280 285
rect 280 284 281 285
rect 281 284 282 285
rect 288 284 289 285
rect 289 284 290 285
rect 290 284 291 285
rect 291 284 292 285
rect 292 284 293 285
rect 337 284 338 285
rect 338 284 339 285
rect 339 284 340 285
rect 340 284 341 285
rect 341 284 342 285
rect 342 284 343 285
rect 343 284 344 285
rect 344 284 345 285
rect 345 284 346 285
rect 346 284 347 285
rect 347 284 348 285
rect 348 284 349 285
rect 349 284 350 285
rect 350 284 351 285
rect 351 284 352 285
rect 361 284 362 285
rect 362 284 363 285
rect 363 284 364 285
rect 364 284 365 285
rect 365 284 366 285
rect 366 284 367 285
rect 377 284 378 285
rect 378 284 379 285
rect 379 284 380 285
rect 380 284 381 285
rect 392 284 393 285
rect 393 284 394 285
rect 394 284 395 285
rect 395 284 396 285
rect 396 284 397 285
rect 397 284 398 285
rect 398 284 399 285
rect 399 284 400 285
rect 400 284 401 285
rect 401 284 402 285
rect 402 284 403 285
rect 403 284 404 285
rect 404 284 405 285
rect 405 284 406 285
rect 50 283 51 284
rect 51 283 52 284
rect 52 283 53 284
rect 53 283 54 284
rect 54 283 55 284
rect 55 283 56 284
rect 56 283 57 284
rect 57 283 58 284
rect 58 283 59 284
rect 163 283 164 284
rect 164 283 165 284
rect 165 283 166 284
rect 166 283 167 284
rect 167 283 168 284
rect 168 283 169 284
rect 169 283 170 284
rect 170 283 171 284
rect 171 283 172 284
rect 173 283 174 284
rect 174 283 175 284
rect 175 283 176 284
rect 176 283 177 284
rect 177 283 178 284
rect 188 283 189 284
rect 189 283 190 284
rect 190 283 191 284
rect 191 283 192 284
rect 192 283 193 284
rect 193 283 194 284
rect 194 283 195 284
rect 195 283 196 284
rect 196 283 197 284
rect 197 283 198 284
rect 238 283 239 284
rect 239 283 240 284
rect 240 283 241 284
rect 241 283 242 284
rect 242 283 243 284
rect 243 283 244 284
rect 244 283 245 284
rect 245 283 246 284
rect 246 283 247 284
rect 247 283 248 284
rect 248 283 249 284
rect 249 283 250 284
rect 250 283 251 284
rect 251 283 252 284
rect 252 283 253 284
rect 253 283 254 284
rect 254 283 255 284
rect 255 283 256 284
rect 256 283 257 284
rect 257 283 258 284
rect 263 283 264 284
rect 264 283 265 284
rect 265 283 266 284
rect 266 283 267 284
rect 267 283 268 284
rect 268 283 269 284
rect 275 283 276 284
rect 276 283 277 284
rect 277 283 278 284
rect 278 283 279 284
rect 279 283 280 284
rect 287 283 288 284
rect 288 283 289 284
rect 289 283 290 284
rect 290 283 291 284
rect 291 283 292 284
rect 292 283 293 284
rect 337 283 338 284
rect 338 283 339 284
rect 339 283 340 284
rect 340 283 341 284
rect 341 283 342 284
rect 342 283 343 284
rect 343 283 344 284
rect 344 283 345 284
rect 345 283 346 284
rect 346 283 347 284
rect 347 283 348 284
rect 348 283 349 284
rect 360 283 361 284
rect 361 283 362 284
rect 362 283 363 284
rect 363 283 364 284
rect 364 283 365 284
rect 365 283 366 284
rect 378 283 379 284
rect 379 283 380 284
rect 380 283 381 284
rect 381 283 382 284
rect 392 283 393 284
rect 393 283 394 284
rect 394 283 395 284
rect 395 283 396 284
rect 396 283 397 284
rect 397 283 398 284
rect 398 283 399 284
rect 399 283 400 284
rect 400 283 401 284
rect 401 283 402 284
rect 402 283 403 284
rect 403 283 404 284
rect 51 282 52 283
rect 52 282 53 283
rect 53 282 54 283
rect 54 282 55 283
rect 55 282 56 283
rect 56 282 57 283
rect 57 282 58 283
rect 58 282 59 283
rect 59 282 60 283
rect 162 282 163 283
rect 163 282 164 283
rect 164 282 165 283
rect 165 282 166 283
rect 166 282 167 283
rect 167 282 168 283
rect 168 282 169 283
rect 169 282 170 283
rect 170 282 171 283
rect 174 282 175 283
rect 175 282 176 283
rect 176 282 177 283
rect 177 282 178 283
rect 190 282 191 283
rect 191 282 192 283
rect 192 282 193 283
rect 193 282 194 283
rect 194 282 195 283
rect 195 282 196 283
rect 196 282 197 283
rect 238 282 239 283
rect 239 282 240 283
rect 240 282 241 283
rect 241 282 242 283
rect 242 282 243 283
rect 243 282 244 283
rect 244 282 245 283
rect 245 282 246 283
rect 246 282 247 283
rect 247 282 248 283
rect 248 282 249 283
rect 249 282 250 283
rect 250 282 251 283
rect 251 282 252 283
rect 252 282 253 283
rect 253 282 254 283
rect 254 282 255 283
rect 263 282 264 283
rect 264 282 265 283
rect 265 282 266 283
rect 266 282 267 283
rect 267 282 268 283
rect 268 282 269 283
rect 269 282 270 283
rect 270 282 271 283
rect 273 282 274 283
rect 274 282 275 283
rect 275 282 276 283
rect 276 282 277 283
rect 277 282 278 283
rect 287 282 288 283
rect 288 282 289 283
rect 289 282 290 283
rect 290 282 291 283
rect 291 282 292 283
rect 292 282 293 283
rect 337 282 338 283
rect 338 282 339 283
rect 339 282 340 283
rect 340 282 341 283
rect 341 282 342 283
rect 342 282 343 283
rect 343 282 344 283
rect 344 282 345 283
rect 345 282 346 283
rect 346 282 347 283
rect 359 282 360 283
rect 360 282 361 283
rect 361 282 362 283
rect 362 282 363 283
rect 363 282 364 283
rect 364 282 365 283
rect 379 282 380 283
rect 380 282 381 283
rect 381 282 382 283
rect 392 282 393 283
rect 393 282 394 283
rect 394 282 395 283
rect 395 282 396 283
rect 396 282 397 283
rect 397 282 398 283
rect 398 282 399 283
rect 399 282 400 283
rect 400 282 401 283
rect 51 281 52 282
rect 52 281 53 282
rect 53 281 54 282
rect 54 281 55 282
rect 55 281 56 282
rect 56 281 57 282
rect 57 281 58 282
rect 58 281 59 282
rect 59 281 60 282
rect 160 281 161 282
rect 161 281 162 282
rect 162 281 163 282
rect 163 281 164 282
rect 164 281 165 282
rect 165 281 166 282
rect 166 281 167 282
rect 167 281 168 282
rect 168 281 169 282
rect 174 281 175 282
rect 175 281 176 282
rect 176 281 177 282
rect 177 281 178 282
rect 178 281 179 282
rect 191 281 192 282
rect 192 281 193 282
rect 193 281 194 282
rect 194 281 195 282
rect 195 281 196 282
rect 241 281 242 282
rect 242 281 243 282
rect 243 281 244 282
rect 244 281 245 282
rect 245 281 246 282
rect 246 281 247 282
rect 247 281 248 282
rect 248 281 249 282
rect 249 281 250 282
rect 250 281 251 282
rect 251 281 252 282
rect 252 281 253 282
rect 253 281 254 282
rect 264 281 265 282
rect 265 281 266 282
rect 266 281 267 282
rect 267 281 268 282
rect 268 281 269 282
rect 269 281 270 282
rect 270 281 271 282
rect 271 281 272 282
rect 272 281 273 282
rect 273 281 274 282
rect 274 281 275 282
rect 275 281 276 282
rect 276 281 277 282
rect 277 281 278 282
rect 287 281 288 282
rect 288 281 289 282
rect 289 281 290 282
rect 290 281 291 282
rect 291 281 292 282
rect 292 281 293 282
rect 338 281 339 282
rect 339 281 340 282
rect 340 281 341 282
rect 341 281 342 282
rect 342 281 343 282
rect 343 281 344 282
rect 344 281 345 282
rect 358 281 359 282
rect 359 281 360 282
rect 360 281 361 282
rect 361 281 362 282
rect 362 281 363 282
rect 363 281 364 282
rect 379 281 380 282
rect 380 281 381 282
rect 381 281 382 282
rect 392 281 393 282
rect 393 281 394 282
rect 394 281 395 282
rect 395 281 396 282
rect 396 281 397 282
rect 397 281 398 282
rect 398 281 399 282
rect 51 280 52 281
rect 52 280 53 281
rect 53 280 54 281
rect 54 280 55 281
rect 55 280 56 281
rect 56 280 57 281
rect 57 280 58 281
rect 58 280 59 281
rect 59 280 60 281
rect 159 280 160 281
rect 160 280 161 281
rect 161 280 162 281
rect 162 280 163 281
rect 163 280 164 281
rect 164 280 165 281
rect 165 280 166 281
rect 166 280 167 281
rect 167 280 168 281
rect 175 280 176 281
rect 176 280 177 281
rect 177 280 178 281
rect 178 280 179 281
rect 179 280 180 281
rect 190 280 191 281
rect 191 280 192 281
rect 192 280 193 281
rect 193 280 194 281
rect 194 280 195 281
rect 249 280 250 281
rect 250 280 251 281
rect 251 280 252 281
rect 252 280 253 281
rect 253 280 254 281
rect 254 280 255 281
rect 265 280 266 281
rect 266 280 267 281
rect 267 280 268 281
rect 268 280 269 281
rect 269 280 270 281
rect 270 280 271 281
rect 271 280 272 281
rect 272 280 273 281
rect 273 280 274 281
rect 274 280 275 281
rect 275 280 276 281
rect 276 280 277 281
rect 277 280 278 281
rect 278 280 279 281
rect 287 280 288 281
rect 288 280 289 281
rect 289 280 290 281
rect 290 280 291 281
rect 291 280 292 281
rect 338 280 339 281
rect 339 280 340 281
rect 340 280 341 281
rect 341 280 342 281
rect 342 280 343 281
rect 358 280 359 281
rect 359 280 360 281
rect 360 280 361 281
rect 361 280 362 281
rect 362 280 363 281
rect 363 280 364 281
rect 380 280 381 281
rect 381 280 382 281
rect 392 280 393 281
rect 393 280 394 281
rect 394 280 395 281
rect 395 280 396 281
rect 396 280 397 281
rect 397 280 398 281
rect 398 280 399 281
rect 51 279 52 280
rect 52 279 53 280
rect 53 279 54 280
rect 54 279 55 280
rect 55 279 56 280
rect 56 279 57 280
rect 57 279 58 280
rect 58 279 59 280
rect 59 279 60 280
rect 60 279 61 280
rect 158 279 159 280
rect 159 279 160 280
rect 160 279 161 280
rect 161 279 162 280
rect 162 279 163 280
rect 163 279 164 280
rect 164 279 165 280
rect 165 279 166 280
rect 175 279 176 280
rect 176 279 177 280
rect 177 279 178 280
rect 178 279 179 280
rect 179 279 180 280
rect 180 279 181 280
rect 189 279 190 280
rect 190 279 191 280
rect 191 279 192 280
rect 192 279 193 280
rect 193 279 194 280
rect 194 279 195 280
rect 249 279 250 280
rect 250 279 251 280
rect 251 279 252 280
rect 252 279 253 280
rect 253 279 254 280
rect 254 279 255 280
rect 265 279 266 280
rect 266 279 267 280
rect 267 279 268 280
rect 268 279 269 280
rect 269 279 270 280
rect 270 279 271 280
rect 271 279 272 280
rect 272 279 273 280
rect 273 279 274 280
rect 274 279 275 280
rect 275 279 276 280
rect 276 279 277 280
rect 277 279 278 280
rect 278 279 279 280
rect 286 279 287 280
rect 287 279 288 280
rect 288 279 289 280
rect 289 279 290 280
rect 290 279 291 280
rect 291 279 292 280
rect 338 279 339 280
rect 339 279 340 280
rect 340 279 341 280
rect 357 279 358 280
rect 358 279 359 280
rect 359 279 360 280
rect 360 279 361 280
rect 361 279 362 280
rect 362 279 363 280
rect 380 279 381 280
rect 381 279 382 280
rect 392 279 393 280
rect 393 279 394 280
rect 394 279 395 280
rect 395 279 396 280
rect 396 279 397 280
rect 397 279 398 280
rect 398 279 399 280
rect 52 278 53 279
rect 53 278 54 279
rect 54 278 55 279
rect 55 278 56 279
rect 56 278 57 279
rect 57 278 58 279
rect 58 278 59 279
rect 59 278 60 279
rect 60 278 61 279
rect 157 278 158 279
rect 158 278 159 279
rect 159 278 160 279
rect 160 278 161 279
rect 161 278 162 279
rect 162 278 163 279
rect 163 278 164 279
rect 164 278 165 279
rect 176 278 177 279
rect 177 278 178 279
rect 178 278 179 279
rect 179 278 180 279
rect 180 278 181 279
rect 181 278 182 279
rect 182 278 183 279
rect 188 278 189 279
rect 189 278 190 279
rect 190 278 191 279
rect 191 278 192 279
rect 192 278 193 279
rect 193 278 194 279
rect 250 278 251 279
rect 251 278 252 279
rect 252 278 253 279
rect 253 278 254 279
rect 254 278 255 279
rect 267 278 268 279
rect 268 278 269 279
rect 269 278 270 279
rect 270 278 271 279
rect 271 278 272 279
rect 272 278 273 279
rect 273 278 274 279
rect 274 278 275 279
rect 275 278 276 279
rect 276 278 277 279
rect 277 278 278 279
rect 286 278 287 279
rect 287 278 288 279
rect 288 278 289 279
rect 289 278 290 279
rect 290 278 291 279
rect 291 278 292 279
rect 338 278 339 279
rect 339 278 340 279
rect 356 278 357 279
rect 357 278 358 279
rect 358 278 359 279
rect 359 278 360 279
rect 360 278 361 279
rect 361 278 362 279
rect 362 278 363 279
rect 381 278 382 279
rect 392 278 393 279
rect 393 278 394 279
rect 394 278 395 279
rect 395 278 396 279
rect 396 278 397 279
rect 397 278 398 279
rect 398 278 399 279
rect 52 277 53 278
rect 53 277 54 278
rect 54 277 55 278
rect 55 277 56 278
rect 56 277 57 278
rect 57 277 58 278
rect 58 277 59 278
rect 59 277 60 278
rect 60 277 61 278
rect 157 277 158 278
rect 158 277 159 278
rect 159 277 160 278
rect 160 277 161 278
rect 161 277 162 278
rect 162 277 163 278
rect 163 277 164 278
rect 177 277 178 278
rect 178 277 179 278
rect 179 277 180 278
rect 180 277 181 278
rect 181 277 182 278
rect 182 277 183 278
rect 183 277 184 278
rect 184 277 185 278
rect 185 277 186 278
rect 186 277 187 278
rect 187 277 188 278
rect 188 277 189 278
rect 189 277 190 278
rect 190 277 191 278
rect 191 277 192 278
rect 192 277 193 278
rect 250 277 251 278
rect 251 277 252 278
rect 252 277 253 278
rect 253 277 254 278
rect 254 277 255 278
rect 255 277 256 278
rect 269 277 270 278
rect 270 277 271 278
rect 271 277 272 278
rect 272 277 273 278
rect 273 277 274 278
rect 274 277 275 278
rect 275 277 276 278
rect 286 277 287 278
rect 287 277 288 278
rect 288 277 289 278
rect 289 277 290 278
rect 290 277 291 278
rect 355 277 356 278
rect 356 277 357 278
rect 357 277 358 278
rect 358 277 359 278
rect 359 277 360 278
rect 360 277 361 278
rect 361 277 362 278
rect 362 277 363 278
rect 381 277 382 278
rect 392 277 393 278
rect 393 277 394 278
rect 394 277 395 278
rect 395 277 396 278
rect 396 277 397 278
rect 397 277 398 278
rect 398 277 399 278
rect 52 276 53 277
rect 53 276 54 277
rect 54 276 55 277
rect 55 276 56 277
rect 56 276 57 277
rect 57 276 58 277
rect 58 276 59 277
rect 59 276 60 277
rect 60 276 61 277
rect 61 276 62 277
rect 156 276 157 277
rect 157 276 158 277
rect 158 276 159 277
rect 159 276 160 277
rect 160 276 161 277
rect 161 276 162 277
rect 162 276 163 277
rect 178 276 179 277
rect 179 276 180 277
rect 180 276 181 277
rect 181 276 182 277
rect 182 276 183 277
rect 183 276 184 277
rect 184 276 185 277
rect 185 276 186 277
rect 186 276 187 277
rect 187 276 188 277
rect 188 276 189 277
rect 189 276 190 277
rect 190 276 191 277
rect 191 276 192 277
rect 250 276 251 277
rect 251 276 252 277
rect 252 276 253 277
rect 253 276 254 277
rect 254 276 255 277
rect 255 276 256 277
rect 285 276 286 277
rect 286 276 287 277
rect 287 276 288 277
rect 288 276 289 277
rect 289 276 290 277
rect 290 276 291 277
rect 354 276 355 277
rect 355 276 356 277
rect 356 276 357 277
rect 357 276 358 277
rect 358 276 359 277
rect 359 276 360 277
rect 360 276 361 277
rect 361 276 362 277
rect 392 276 393 277
rect 393 276 394 277
rect 394 276 395 277
rect 395 276 396 277
rect 396 276 397 277
rect 397 276 398 277
rect 53 275 54 276
rect 54 275 55 276
rect 55 275 56 276
rect 56 275 57 276
rect 57 275 58 276
rect 58 275 59 276
rect 59 275 60 276
rect 60 275 61 276
rect 61 275 62 276
rect 155 275 156 276
rect 156 275 157 276
rect 157 275 158 276
rect 158 275 159 276
rect 159 275 160 276
rect 160 275 161 276
rect 161 275 162 276
rect 180 275 181 276
rect 181 275 182 276
rect 182 275 183 276
rect 183 275 184 276
rect 184 275 185 276
rect 185 275 186 276
rect 186 275 187 276
rect 187 275 188 276
rect 188 275 189 276
rect 189 275 190 276
rect 190 275 191 276
rect 251 275 252 276
rect 252 275 253 276
rect 253 275 254 276
rect 254 275 255 276
rect 255 275 256 276
rect 256 275 257 276
rect 284 275 285 276
rect 285 275 286 276
rect 286 275 287 276
rect 287 275 288 276
rect 288 275 289 276
rect 289 275 290 276
rect 353 275 354 276
rect 354 275 355 276
rect 355 275 356 276
rect 356 275 357 276
rect 357 275 358 276
rect 358 275 359 276
rect 359 275 360 276
rect 360 275 361 276
rect 361 275 362 276
rect 391 275 392 276
rect 392 275 393 276
rect 393 275 394 276
rect 394 275 395 276
rect 395 275 396 276
rect 396 275 397 276
rect 397 275 398 276
rect 53 274 54 275
rect 54 274 55 275
rect 55 274 56 275
rect 56 274 57 275
rect 57 274 58 275
rect 58 274 59 275
rect 59 274 60 275
rect 60 274 61 275
rect 61 274 62 275
rect 155 274 156 275
rect 156 274 157 275
rect 157 274 158 275
rect 158 274 159 275
rect 159 274 160 275
rect 160 274 161 275
rect 182 274 183 275
rect 183 274 184 275
rect 184 274 185 275
rect 185 274 186 275
rect 186 274 187 275
rect 187 274 188 275
rect 188 274 189 275
rect 189 274 190 275
rect 190 274 191 275
rect 251 274 252 275
rect 252 274 253 275
rect 253 274 254 275
rect 254 274 255 275
rect 255 274 256 275
rect 256 274 257 275
rect 257 274 258 275
rect 283 274 284 275
rect 284 274 285 275
rect 285 274 286 275
rect 286 274 287 275
rect 287 274 288 275
rect 288 274 289 275
rect 289 274 290 275
rect 353 274 354 275
rect 354 274 355 275
rect 355 274 356 275
rect 356 274 357 275
rect 357 274 358 275
rect 358 274 359 275
rect 359 274 360 275
rect 360 274 361 275
rect 361 274 362 275
rect 362 274 363 275
rect 391 274 392 275
rect 392 274 393 275
rect 393 274 394 275
rect 394 274 395 275
rect 395 274 396 275
rect 396 274 397 275
rect 397 274 398 275
rect 53 273 54 274
rect 54 273 55 274
rect 55 273 56 274
rect 56 273 57 274
rect 57 273 58 274
rect 58 273 59 274
rect 59 273 60 274
rect 60 273 61 274
rect 61 273 62 274
rect 62 273 63 274
rect 154 273 155 274
rect 155 273 156 274
rect 156 273 157 274
rect 157 273 158 274
rect 158 273 159 274
rect 159 273 160 274
rect 160 273 161 274
rect 185 273 186 274
rect 186 273 187 274
rect 187 273 188 274
rect 188 273 189 274
rect 189 273 190 274
rect 252 273 253 274
rect 253 273 254 274
rect 254 273 255 274
rect 255 273 256 274
rect 256 273 257 274
rect 257 273 258 274
rect 258 273 259 274
rect 283 273 284 274
rect 284 273 285 274
rect 285 273 286 274
rect 286 273 287 274
rect 287 273 288 274
rect 288 273 289 274
rect 352 273 353 274
rect 353 273 354 274
rect 354 273 355 274
rect 355 273 356 274
rect 356 273 357 274
rect 357 273 358 274
rect 358 273 359 274
rect 359 273 360 274
rect 360 273 361 274
rect 361 273 362 274
rect 362 273 363 274
rect 391 273 392 274
rect 392 273 393 274
rect 393 273 394 274
rect 394 273 395 274
rect 395 273 396 274
rect 396 273 397 274
rect 397 273 398 274
rect 54 272 55 273
rect 55 272 56 273
rect 56 272 57 273
rect 57 272 58 273
rect 58 272 59 273
rect 59 272 60 273
rect 60 272 61 273
rect 61 272 62 273
rect 62 272 63 273
rect 154 272 155 273
rect 155 272 156 273
rect 156 272 157 273
rect 157 272 158 273
rect 158 272 159 273
rect 159 272 160 273
rect 184 272 185 273
rect 185 272 186 273
rect 186 272 187 273
rect 187 272 188 273
rect 188 272 189 273
rect 189 272 190 273
rect 253 272 254 273
rect 254 272 255 273
rect 255 272 256 273
rect 256 272 257 273
rect 257 272 258 273
rect 258 272 259 273
rect 259 272 260 273
rect 281 272 282 273
rect 282 272 283 273
rect 283 272 284 273
rect 284 272 285 273
rect 285 272 286 273
rect 286 272 287 273
rect 287 272 288 273
rect 288 272 289 273
rect 351 272 352 273
rect 352 272 353 273
rect 357 272 358 273
rect 358 272 359 273
rect 359 272 360 273
rect 360 272 361 273
rect 361 272 362 273
rect 362 272 363 273
rect 363 272 364 273
rect 391 272 392 273
rect 392 272 393 273
rect 393 272 394 273
rect 394 272 395 273
rect 395 272 396 273
rect 396 272 397 273
rect 397 272 398 273
rect 54 271 55 272
rect 55 271 56 272
rect 56 271 57 272
rect 57 271 58 272
rect 58 271 59 272
rect 59 271 60 272
rect 60 271 61 272
rect 61 271 62 272
rect 62 271 63 272
rect 63 271 64 272
rect 153 271 154 272
rect 154 271 155 272
rect 155 271 156 272
rect 156 271 157 272
rect 157 271 158 272
rect 158 271 159 272
rect 184 271 185 272
rect 185 271 186 272
rect 186 271 187 272
rect 187 271 188 272
rect 188 271 189 272
rect 253 271 254 272
rect 254 271 255 272
rect 255 271 256 272
rect 256 271 257 272
rect 257 271 258 272
rect 258 271 259 272
rect 259 271 260 272
rect 260 271 261 272
rect 280 271 281 272
rect 281 271 282 272
rect 282 271 283 272
rect 283 271 284 272
rect 284 271 285 272
rect 285 271 286 272
rect 286 271 287 272
rect 287 271 288 272
rect 351 271 352 272
rect 358 271 359 272
rect 359 271 360 272
rect 360 271 361 272
rect 361 271 362 272
rect 362 271 363 272
rect 363 271 364 272
rect 364 271 365 272
rect 390 271 391 272
rect 391 271 392 272
rect 392 271 393 272
rect 393 271 394 272
rect 394 271 395 272
rect 395 271 396 272
rect 396 271 397 272
rect 55 270 56 271
rect 56 270 57 271
rect 57 270 58 271
rect 58 270 59 271
rect 59 270 60 271
rect 60 270 61 271
rect 61 270 62 271
rect 62 270 63 271
rect 63 270 64 271
rect 153 270 154 271
rect 154 270 155 271
rect 155 270 156 271
rect 156 270 157 271
rect 157 270 158 271
rect 158 270 159 271
rect 183 270 184 271
rect 184 270 185 271
rect 185 270 186 271
rect 186 270 187 271
rect 187 270 188 271
rect 188 270 189 271
rect 254 270 255 271
rect 255 270 256 271
rect 256 270 257 271
rect 257 270 258 271
rect 258 270 259 271
rect 259 270 260 271
rect 260 270 261 271
rect 261 270 262 271
rect 262 270 263 271
rect 278 270 279 271
rect 279 270 280 271
rect 280 270 281 271
rect 281 270 282 271
rect 282 270 283 271
rect 283 270 284 271
rect 284 270 285 271
rect 285 270 286 271
rect 286 270 287 271
rect 359 270 360 271
rect 360 270 361 271
rect 361 270 362 271
rect 362 270 363 271
rect 363 270 364 271
rect 364 270 365 271
rect 365 270 366 271
rect 366 270 367 271
rect 390 270 391 271
rect 391 270 392 271
rect 392 270 393 271
rect 393 270 394 271
rect 394 270 395 271
rect 395 270 396 271
rect 396 270 397 271
rect 55 269 56 270
rect 56 269 57 270
rect 57 269 58 270
rect 58 269 59 270
rect 59 269 60 270
rect 60 269 61 270
rect 61 269 62 270
rect 62 269 63 270
rect 63 269 64 270
rect 64 269 65 270
rect 152 269 153 270
rect 153 269 154 270
rect 154 269 155 270
rect 155 269 156 270
rect 156 269 157 270
rect 157 269 158 270
rect 183 269 184 270
rect 184 269 185 270
rect 185 269 186 270
rect 186 269 187 270
rect 187 269 188 270
rect 188 269 189 270
rect 255 269 256 270
rect 256 269 257 270
rect 257 269 258 270
rect 258 269 259 270
rect 259 269 260 270
rect 260 269 261 270
rect 261 269 262 270
rect 262 269 263 270
rect 263 269 264 270
rect 264 269 265 270
rect 276 269 277 270
rect 277 269 278 270
rect 278 269 279 270
rect 279 269 280 270
rect 280 269 281 270
rect 281 269 282 270
rect 282 269 283 270
rect 283 269 284 270
rect 284 269 285 270
rect 285 269 286 270
rect 359 269 360 270
rect 360 269 361 270
rect 361 269 362 270
rect 362 269 363 270
rect 363 269 364 270
rect 364 269 365 270
rect 365 269 366 270
rect 366 269 367 270
rect 367 269 368 270
rect 368 269 369 270
rect 390 269 391 270
rect 391 269 392 270
rect 392 269 393 270
rect 393 269 394 270
rect 394 269 395 270
rect 395 269 396 270
rect 396 269 397 270
rect 55 268 56 269
rect 56 268 57 269
rect 57 268 58 269
rect 58 268 59 269
rect 59 268 60 269
rect 60 268 61 269
rect 61 268 62 269
rect 62 268 63 269
rect 63 268 64 269
rect 64 268 65 269
rect 152 268 153 269
rect 153 268 154 269
rect 154 268 155 269
rect 155 268 156 269
rect 156 268 157 269
rect 157 268 158 269
rect 182 268 183 269
rect 183 268 184 269
rect 184 268 185 269
rect 185 268 186 269
rect 186 268 187 269
rect 187 268 188 269
rect 256 268 257 269
rect 257 268 258 269
rect 258 268 259 269
rect 259 268 260 269
rect 260 268 261 269
rect 261 268 262 269
rect 262 268 263 269
rect 263 268 264 269
rect 264 268 265 269
rect 265 268 266 269
rect 266 268 267 269
rect 267 268 268 269
rect 268 268 269 269
rect 269 268 270 269
rect 270 268 271 269
rect 271 268 272 269
rect 272 268 273 269
rect 273 268 274 269
rect 274 268 275 269
rect 275 268 276 269
rect 276 268 277 269
rect 277 268 278 269
rect 278 268 279 269
rect 279 268 280 269
rect 280 268 281 269
rect 281 268 282 269
rect 282 268 283 269
rect 283 268 284 269
rect 284 268 285 269
rect 359 268 360 269
rect 360 268 361 269
rect 361 268 362 269
rect 362 268 363 269
rect 363 268 364 269
rect 364 268 365 269
rect 365 268 366 269
rect 366 268 367 269
rect 367 268 368 269
rect 368 268 369 269
rect 369 268 370 269
rect 389 268 390 269
rect 390 268 391 269
rect 391 268 392 269
rect 392 268 393 269
rect 393 268 394 269
rect 394 268 395 269
rect 395 268 396 269
rect 56 267 57 268
rect 57 267 58 268
rect 58 267 59 268
rect 59 267 60 268
rect 60 267 61 268
rect 61 267 62 268
rect 62 267 63 268
rect 63 267 64 268
rect 64 267 65 268
rect 65 267 66 268
rect 151 267 152 268
rect 152 267 153 268
rect 153 267 154 268
rect 154 267 155 268
rect 155 267 156 268
rect 156 267 157 268
rect 182 267 183 268
rect 183 267 184 268
rect 184 267 185 268
rect 185 267 186 268
rect 186 267 187 268
rect 187 267 188 268
rect 258 267 259 268
rect 259 267 260 268
rect 260 267 261 268
rect 261 267 262 268
rect 262 267 263 268
rect 263 267 264 268
rect 264 267 265 268
rect 265 267 266 268
rect 266 267 267 268
rect 267 267 268 268
rect 268 267 269 268
rect 269 267 270 268
rect 270 267 271 268
rect 271 267 272 268
rect 272 267 273 268
rect 273 267 274 268
rect 274 267 275 268
rect 275 267 276 268
rect 276 267 277 268
rect 277 267 278 268
rect 278 267 279 268
rect 279 267 280 268
rect 280 267 281 268
rect 281 267 282 268
rect 282 267 283 268
rect 283 267 284 268
rect 359 267 360 268
rect 360 267 361 268
rect 361 267 362 268
rect 362 267 363 268
rect 363 267 364 268
rect 364 267 365 268
rect 365 267 366 268
rect 366 267 367 268
rect 367 267 368 268
rect 368 267 369 268
rect 369 267 370 268
rect 370 267 371 268
rect 389 267 390 268
rect 390 267 391 268
rect 391 267 392 268
rect 392 267 393 268
rect 393 267 394 268
rect 394 267 395 268
rect 395 267 396 268
rect 56 266 57 267
rect 57 266 58 267
rect 58 266 59 267
rect 59 266 60 267
rect 60 266 61 267
rect 61 266 62 267
rect 62 266 63 267
rect 63 266 64 267
rect 64 266 65 267
rect 65 266 66 267
rect 151 266 152 267
rect 152 266 153 267
rect 153 266 154 267
rect 154 266 155 267
rect 155 266 156 267
rect 156 266 157 267
rect 173 266 174 267
rect 174 266 175 267
rect 175 266 176 267
rect 176 266 177 267
rect 177 266 178 267
rect 178 266 179 267
rect 179 266 180 267
rect 180 266 181 267
rect 181 266 182 267
rect 182 266 183 267
rect 183 266 184 267
rect 184 266 185 267
rect 185 266 186 267
rect 186 266 187 267
rect 187 266 188 267
rect 225 266 226 267
rect 226 266 227 267
rect 227 266 228 267
rect 228 266 229 267
rect 229 266 230 267
rect 230 266 231 267
rect 231 266 232 267
rect 232 266 233 267
rect 259 266 260 267
rect 260 266 261 267
rect 261 266 262 267
rect 262 266 263 267
rect 263 266 264 267
rect 264 266 265 267
rect 265 266 266 267
rect 266 266 267 267
rect 267 266 268 267
rect 268 266 269 267
rect 269 266 270 267
rect 270 266 271 267
rect 271 266 272 267
rect 272 266 273 267
rect 273 266 274 267
rect 274 266 275 267
rect 275 266 276 267
rect 276 266 277 267
rect 277 266 278 267
rect 278 266 279 267
rect 279 266 280 267
rect 280 266 281 267
rect 281 266 282 267
rect 359 266 360 267
rect 360 266 361 267
rect 361 266 362 267
rect 362 266 363 267
rect 363 266 364 267
rect 364 266 365 267
rect 365 266 366 267
rect 366 266 367 267
rect 367 266 368 267
rect 368 266 369 267
rect 369 266 370 267
rect 370 266 371 267
rect 371 266 372 267
rect 389 266 390 267
rect 390 266 391 267
rect 391 266 392 267
rect 392 266 393 267
rect 393 266 394 267
rect 394 266 395 267
rect 395 266 396 267
rect 57 265 58 266
rect 58 265 59 266
rect 59 265 60 266
rect 60 265 61 266
rect 61 265 62 266
rect 62 265 63 266
rect 63 265 64 266
rect 64 265 65 266
rect 65 265 66 266
rect 66 265 67 266
rect 151 265 152 266
rect 152 265 153 266
rect 153 265 154 266
rect 154 265 155 266
rect 155 265 156 266
rect 156 265 157 266
rect 169 265 170 266
rect 170 265 171 266
rect 171 265 172 266
rect 172 265 173 266
rect 173 265 174 266
rect 174 265 175 266
rect 175 265 176 266
rect 176 265 177 266
rect 177 265 178 266
rect 178 265 179 266
rect 179 265 180 266
rect 180 265 181 266
rect 181 265 182 266
rect 182 265 183 266
rect 183 265 184 266
rect 184 265 185 266
rect 185 265 186 266
rect 186 265 187 266
rect 187 265 188 266
rect 225 265 226 266
rect 226 265 227 266
rect 227 265 228 266
rect 228 265 229 266
rect 229 265 230 266
rect 230 265 231 266
rect 231 265 232 266
rect 232 265 233 266
rect 233 265 234 266
rect 234 265 235 266
rect 235 265 236 266
rect 261 265 262 266
rect 262 265 263 266
rect 263 265 264 266
rect 264 265 265 266
rect 265 265 266 266
rect 266 265 267 266
rect 267 265 268 266
rect 268 265 269 266
rect 269 265 270 266
rect 270 265 271 266
rect 271 265 272 266
rect 272 265 273 266
rect 273 265 274 266
rect 274 265 275 266
rect 275 265 276 266
rect 276 265 277 266
rect 277 265 278 266
rect 278 265 279 266
rect 279 265 280 266
rect 359 265 360 266
rect 360 265 361 266
rect 361 265 362 266
rect 362 265 363 266
rect 363 265 364 266
rect 364 265 365 266
rect 365 265 366 266
rect 366 265 367 266
rect 367 265 368 266
rect 368 265 369 266
rect 369 265 370 266
rect 370 265 371 266
rect 371 265 372 266
rect 372 265 373 266
rect 388 265 389 266
rect 389 265 390 266
rect 390 265 391 266
rect 391 265 392 266
rect 392 265 393 266
rect 393 265 394 266
rect 394 265 395 266
rect 57 264 58 265
rect 58 264 59 265
rect 59 264 60 265
rect 60 264 61 265
rect 61 264 62 265
rect 62 264 63 265
rect 63 264 64 265
rect 64 264 65 265
rect 65 264 66 265
rect 66 264 67 265
rect 150 264 151 265
rect 151 264 152 265
rect 152 264 153 265
rect 153 264 154 265
rect 154 264 155 265
rect 155 264 156 265
rect 156 264 157 265
rect 165 264 166 265
rect 166 264 167 265
rect 167 264 168 265
rect 168 264 169 265
rect 169 264 170 265
rect 170 264 171 265
rect 171 264 172 265
rect 172 264 173 265
rect 173 264 174 265
rect 174 264 175 265
rect 175 264 176 265
rect 176 264 177 265
rect 177 264 178 265
rect 178 264 179 265
rect 179 264 180 265
rect 180 264 181 265
rect 181 264 182 265
rect 182 264 183 265
rect 183 264 184 265
rect 184 264 185 265
rect 185 264 186 265
rect 186 264 187 265
rect 224 264 225 265
rect 225 264 226 265
rect 226 264 227 265
rect 227 264 228 265
rect 228 264 229 265
rect 229 264 230 265
rect 230 264 231 265
rect 231 264 232 265
rect 232 264 233 265
rect 233 264 234 265
rect 234 264 235 265
rect 235 264 236 265
rect 236 264 237 265
rect 237 264 238 265
rect 263 264 264 265
rect 264 264 265 265
rect 265 264 266 265
rect 266 264 267 265
rect 267 264 268 265
rect 268 264 269 265
rect 269 264 270 265
rect 270 264 271 265
rect 271 264 272 265
rect 272 264 273 265
rect 273 264 274 265
rect 274 264 275 265
rect 275 264 276 265
rect 276 264 277 265
rect 277 264 278 265
rect 358 264 359 265
rect 359 264 360 265
rect 360 264 361 265
rect 361 264 362 265
rect 362 264 363 265
rect 363 264 364 265
rect 364 264 365 265
rect 369 264 370 265
rect 370 264 371 265
rect 371 264 372 265
rect 372 264 373 265
rect 388 264 389 265
rect 389 264 390 265
rect 390 264 391 265
rect 391 264 392 265
rect 392 264 393 265
rect 393 264 394 265
rect 394 264 395 265
rect 58 263 59 264
rect 59 263 60 264
rect 60 263 61 264
rect 61 263 62 264
rect 62 263 63 264
rect 63 263 64 264
rect 64 263 65 264
rect 65 263 66 264
rect 66 263 67 264
rect 67 263 68 264
rect 150 263 151 264
rect 151 263 152 264
rect 152 263 153 264
rect 153 263 154 264
rect 154 263 155 264
rect 155 263 156 264
rect 162 263 163 264
rect 163 263 164 264
rect 164 263 165 264
rect 165 263 166 264
rect 166 263 167 264
rect 167 263 168 264
rect 168 263 169 264
rect 169 263 170 264
rect 170 263 171 264
rect 171 263 172 264
rect 172 263 173 264
rect 173 263 174 264
rect 174 263 175 264
rect 175 263 176 264
rect 176 263 177 264
rect 177 263 178 264
rect 178 263 179 264
rect 179 263 180 264
rect 180 263 181 264
rect 181 263 182 264
rect 182 263 183 264
rect 183 263 184 264
rect 184 263 185 264
rect 185 263 186 264
rect 186 263 187 264
rect 226 263 227 264
rect 227 263 228 264
rect 228 263 229 264
rect 229 263 230 264
rect 230 263 231 264
rect 231 263 232 264
rect 232 263 233 264
rect 233 263 234 264
rect 234 263 235 264
rect 235 263 236 264
rect 236 263 237 264
rect 237 263 238 264
rect 238 263 239 264
rect 239 263 240 264
rect 267 263 268 264
rect 268 263 269 264
rect 269 263 270 264
rect 270 263 271 264
rect 271 263 272 264
rect 272 263 273 264
rect 273 263 274 264
rect 358 263 359 264
rect 359 263 360 264
rect 360 263 361 264
rect 361 263 362 264
rect 362 263 363 264
rect 363 263 364 264
rect 371 263 372 264
rect 387 263 388 264
rect 388 263 389 264
rect 389 263 390 264
rect 390 263 391 264
rect 391 263 392 264
rect 392 263 393 264
rect 393 263 394 264
rect 58 262 59 263
rect 59 262 60 263
rect 60 262 61 263
rect 61 262 62 263
rect 62 262 63 263
rect 63 262 64 263
rect 64 262 65 263
rect 65 262 66 263
rect 66 262 67 263
rect 67 262 68 263
rect 68 262 69 263
rect 110 262 111 263
rect 111 262 112 263
rect 150 262 151 263
rect 151 262 152 263
rect 152 262 153 263
rect 153 262 154 263
rect 154 262 155 263
rect 155 262 156 263
rect 160 262 161 263
rect 161 262 162 263
rect 162 262 163 263
rect 163 262 164 263
rect 164 262 165 263
rect 165 262 166 263
rect 166 262 167 263
rect 167 262 168 263
rect 168 262 169 263
rect 169 262 170 263
rect 170 262 171 263
rect 171 262 172 263
rect 172 262 173 263
rect 173 262 174 263
rect 174 262 175 263
rect 175 262 176 263
rect 176 262 177 263
rect 177 262 178 263
rect 178 262 179 263
rect 179 262 180 263
rect 180 262 181 263
rect 181 262 182 263
rect 182 262 183 263
rect 183 262 184 263
rect 184 262 185 263
rect 185 262 186 263
rect 186 262 187 263
rect 227 262 228 263
rect 228 262 229 263
rect 229 262 230 263
rect 230 262 231 263
rect 231 262 232 263
rect 232 262 233 263
rect 237 262 238 263
rect 238 262 239 263
rect 239 262 240 263
rect 240 262 241 263
rect 357 262 358 263
rect 358 262 359 263
rect 359 262 360 263
rect 360 262 361 263
rect 361 262 362 263
rect 362 262 363 263
rect 387 262 388 263
rect 388 262 389 263
rect 389 262 390 263
rect 390 262 391 263
rect 391 262 392 263
rect 392 262 393 263
rect 393 262 394 263
rect 59 261 60 262
rect 60 261 61 262
rect 61 261 62 262
rect 62 261 63 262
rect 63 261 64 262
rect 64 261 65 262
rect 65 261 66 262
rect 66 261 67 262
rect 67 261 68 262
rect 68 261 69 262
rect 110 261 111 262
rect 111 261 112 262
rect 112 261 113 262
rect 113 261 114 262
rect 149 261 150 262
rect 150 261 151 262
rect 151 261 152 262
rect 152 261 153 262
rect 153 261 154 262
rect 154 261 155 262
rect 155 261 156 262
rect 156 261 157 262
rect 157 261 158 262
rect 158 261 159 262
rect 159 261 160 262
rect 160 261 161 262
rect 161 261 162 262
rect 162 261 163 262
rect 163 261 164 262
rect 164 261 165 262
rect 165 261 166 262
rect 166 261 167 262
rect 167 261 168 262
rect 168 261 169 262
rect 169 261 170 262
rect 170 261 171 262
rect 171 261 172 262
rect 172 261 173 262
rect 173 261 174 262
rect 174 261 175 262
rect 175 261 176 262
rect 176 261 177 262
rect 177 261 178 262
rect 178 261 179 262
rect 179 261 180 262
rect 180 261 181 262
rect 181 261 182 262
rect 182 261 183 262
rect 183 261 184 262
rect 184 261 185 262
rect 185 261 186 262
rect 186 261 187 262
rect 228 261 229 262
rect 229 261 230 262
rect 230 261 231 262
rect 231 261 232 262
rect 240 261 241 262
rect 241 261 242 262
rect 346 261 347 262
rect 355 261 356 262
rect 356 261 357 262
rect 357 261 358 262
rect 358 261 359 262
rect 359 261 360 262
rect 360 261 361 262
rect 361 261 362 262
rect 362 261 363 262
rect 386 261 387 262
rect 387 261 388 262
rect 388 261 389 262
rect 389 261 390 262
rect 390 261 391 262
rect 391 261 392 262
rect 392 261 393 262
rect 59 260 60 261
rect 60 260 61 261
rect 61 260 62 261
rect 62 260 63 261
rect 63 260 64 261
rect 64 260 65 261
rect 65 260 66 261
rect 66 260 67 261
rect 67 260 68 261
rect 68 260 69 261
rect 69 260 70 261
rect 111 260 112 261
rect 112 260 113 261
rect 113 260 114 261
rect 114 260 115 261
rect 149 260 150 261
rect 150 260 151 261
rect 151 260 152 261
rect 152 260 153 261
rect 153 260 154 261
rect 154 260 155 261
rect 155 260 156 261
rect 156 260 157 261
rect 157 260 158 261
rect 158 260 159 261
rect 159 260 160 261
rect 160 260 161 261
rect 161 260 162 261
rect 162 260 163 261
rect 163 260 164 261
rect 164 260 165 261
rect 165 260 166 261
rect 166 260 167 261
rect 167 260 168 261
rect 168 260 169 261
rect 169 260 170 261
rect 170 260 171 261
rect 171 260 172 261
rect 172 260 173 261
rect 173 260 174 261
rect 174 260 175 261
rect 175 260 176 261
rect 176 260 177 261
rect 177 260 178 261
rect 178 260 179 261
rect 179 260 180 261
rect 180 260 181 261
rect 181 260 182 261
rect 182 260 183 261
rect 183 260 184 261
rect 184 260 185 261
rect 185 260 186 261
rect 186 260 187 261
rect 228 260 229 261
rect 229 260 230 261
rect 230 260 231 261
rect 231 260 232 261
rect 232 260 233 261
rect 316 260 317 261
rect 345 260 346 261
rect 346 260 347 261
rect 347 260 348 261
rect 348 260 349 261
rect 349 260 350 261
rect 350 260 351 261
rect 352 260 353 261
rect 353 260 354 261
rect 354 260 355 261
rect 355 260 356 261
rect 356 260 357 261
rect 357 260 358 261
rect 358 260 359 261
rect 359 260 360 261
rect 360 260 361 261
rect 361 260 362 261
rect 386 260 387 261
rect 387 260 388 261
rect 388 260 389 261
rect 389 260 390 261
rect 390 260 391 261
rect 391 260 392 261
rect 392 260 393 261
rect 60 259 61 260
rect 61 259 62 260
rect 62 259 63 260
rect 63 259 64 260
rect 64 259 65 260
rect 65 259 66 260
rect 66 259 67 260
rect 67 259 68 260
rect 68 259 69 260
rect 69 259 70 260
rect 70 259 71 260
rect 111 259 112 260
rect 112 259 113 260
rect 113 259 114 260
rect 114 259 115 260
rect 115 259 116 260
rect 116 259 117 260
rect 117 259 118 260
rect 149 259 150 260
rect 150 259 151 260
rect 151 259 152 260
rect 152 259 153 260
rect 153 259 154 260
rect 154 259 155 260
rect 155 259 156 260
rect 156 259 157 260
rect 157 259 158 260
rect 158 259 159 260
rect 159 259 160 260
rect 160 259 161 260
rect 161 259 162 260
rect 162 259 163 260
rect 163 259 164 260
rect 164 259 165 260
rect 165 259 166 260
rect 166 259 167 260
rect 167 259 168 260
rect 168 259 169 260
rect 169 259 170 260
rect 175 259 176 260
rect 176 259 177 260
rect 177 259 178 260
rect 178 259 179 260
rect 179 259 180 260
rect 180 259 181 260
rect 181 259 182 260
rect 182 259 183 260
rect 183 259 184 260
rect 184 259 185 260
rect 185 259 186 260
rect 186 259 187 260
rect 228 259 229 260
rect 229 259 230 260
rect 230 259 231 260
rect 231 259 232 260
rect 232 259 233 260
rect 233 259 234 260
rect 234 259 235 260
rect 235 259 236 260
rect 236 259 237 260
rect 237 259 238 260
rect 238 259 239 260
rect 316 259 317 260
rect 345 259 346 260
rect 346 259 347 260
rect 347 259 348 260
rect 348 259 349 260
rect 349 259 350 260
rect 350 259 351 260
rect 351 259 352 260
rect 352 259 353 260
rect 353 259 354 260
rect 354 259 355 260
rect 355 259 356 260
rect 356 259 357 260
rect 357 259 358 260
rect 358 259 359 260
rect 359 259 360 260
rect 360 259 361 260
rect 385 259 386 260
rect 386 259 387 260
rect 387 259 388 260
rect 388 259 389 260
rect 389 259 390 260
rect 390 259 391 260
rect 391 259 392 260
rect 61 258 62 259
rect 62 258 63 259
rect 63 258 64 259
rect 64 258 65 259
rect 65 258 66 259
rect 66 258 67 259
rect 67 258 68 259
rect 68 258 69 259
rect 69 258 70 259
rect 70 258 71 259
rect 112 258 113 259
rect 113 258 114 259
rect 114 258 115 259
rect 115 258 116 259
rect 116 258 117 259
rect 117 258 118 259
rect 118 258 119 259
rect 119 258 120 259
rect 120 258 121 259
rect 146 258 147 259
rect 147 258 148 259
rect 148 258 149 259
rect 149 258 150 259
rect 150 258 151 259
rect 151 258 152 259
rect 152 258 153 259
rect 153 258 154 259
rect 154 258 155 259
rect 155 258 156 259
rect 156 258 157 259
rect 157 258 158 259
rect 158 258 159 259
rect 159 258 160 259
rect 160 258 161 259
rect 161 258 162 259
rect 162 258 163 259
rect 163 258 164 259
rect 178 258 179 259
rect 179 258 180 259
rect 180 258 181 259
rect 181 258 182 259
rect 182 258 183 259
rect 183 258 184 259
rect 184 258 185 259
rect 185 258 186 259
rect 186 258 187 259
rect 228 258 229 259
rect 229 258 230 259
rect 230 258 231 259
rect 231 258 232 259
rect 232 258 233 259
rect 233 258 234 259
rect 234 258 235 259
rect 235 258 236 259
rect 236 258 237 259
rect 237 258 238 259
rect 238 258 239 259
rect 239 258 240 259
rect 240 258 241 259
rect 241 258 242 259
rect 316 258 317 259
rect 346 258 347 259
rect 347 258 348 259
rect 348 258 349 259
rect 349 258 350 259
rect 350 258 351 259
rect 351 258 352 259
rect 352 258 353 259
rect 353 258 354 259
rect 354 258 355 259
rect 355 258 356 259
rect 356 258 357 259
rect 357 258 358 259
rect 358 258 359 259
rect 359 258 360 259
rect 385 258 386 259
rect 386 258 387 259
rect 387 258 388 259
rect 388 258 389 259
rect 389 258 390 259
rect 390 258 391 259
rect 391 258 392 259
rect 61 257 62 258
rect 62 257 63 258
rect 63 257 64 258
rect 64 257 65 258
rect 65 257 66 258
rect 66 257 67 258
rect 67 257 68 258
rect 68 257 69 258
rect 69 257 70 258
rect 70 257 71 258
rect 71 257 72 258
rect 112 257 113 258
rect 113 257 114 258
rect 114 257 115 258
rect 115 257 116 258
rect 116 257 117 258
rect 117 257 118 258
rect 118 257 119 258
rect 119 257 120 258
rect 120 257 121 258
rect 121 257 122 258
rect 122 257 123 258
rect 123 257 124 258
rect 141 257 142 258
rect 142 257 143 258
rect 143 257 144 258
rect 144 257 145 258
rect 145 257 146 258
rect 146 257 147 258
rect 147 257 148 258
rect 148 257 149 258
rect 149 257 150 258
rect 150 257 151 258
rect 151 257 152 258
rect 152 257 153 258
rect 153 257 154 258
rect 154 257 155 258
rect 155 257 156 258
rect 156 257 157 258
rect 157 257 158 258
rect 158 257 159 258
rect 159 257 160 258
rect 170 257 171 258
rect 171 257 172 258
rect 172 257 173 258
rect 173 257 174 258
rect 174 257 175 258
rect 175 257 176 258
rect 176 257 177 258
rect 177 257 178 258
rect 178 257 179 258
rect 179 257 180 258
rect 180 257 181 258
rect 181 257 182 258
rect 182 257 183 258
rect 183 257 184 258
rect 184 257 185 258
rect 185 257 186 258
rect 186 257 187 258
rect 228 257 229 258
rect 229 257 230 258
rect 230 257 231 258
rect 231 257 232 258
rect 232 257 233 258
rect 233 257 234 258
rect 234 257 235 258
rect 235 257 236 258
rect 236 257 237 258
rect 237 257 238 258
rect 238 257 239 258
rect 239 257 240 258
rect 240 257 241 258
rect 241 257 242 258
rect 242 257 243 258
rect 243 257 244 258
rect 316 257 317 258
rect 317 257 318 258
rect 347 257 348 258
rect 348 257 349 258
rect 349 257 350 258
rect 350 257 351 258
rect 351 257 352 258
rect 352 257 353 258
rect 353 257 354 258
rect 354 257 355 258
rect 355 257 356 258
rect 356 257 357 258
rect 357 257 358 258
rect 358 257 359 258
rect 384 257 385 258
rect 385 257 386 258
rect 386 257 387 258
rect 387 257 388 258
rect 388 257 389 258
rect 389 257 390 258
rect 390 257 391 258
rect 62 256 63 257
rect 63 256 64 257
rect 64 256 65 257
rect 65 256 66 257
rect 66 256 67 257
rect 67 256 68 257
rect 68 256 69 257
rect 69 256 70 257
rect 70 256 71 257
rect 71 256 72 257
rect 72 256 73 257
rect 112 256 113 257
rect 113 256 114 257
rect 114 256 115 257
rect 115 256 116 257
rect 116 256 117 257
rect 117 256 118 257
rect 118 256 119 257
rect 119 256 120 257
rect 120 256 121 257
rect 121 256 122 257
rect 122 256 123 257
rect 123 256 124 257
rect 124 256 125 257
rect 125 256 126 257
rect 126 256 127 257
rect 127 256 128 257
rect 128 256 129 257
rect 129 256 130 257
rect 130 256 131 257
rect 131 256 132 257
rect 132 256 133 257
rect 133 256 134 257
rect 134 256 135 257
rect 135 256 136 257
rect 136 256 137 257
rect 137 256 138 257
rect 138 256 139 257
rect 139 256 140 257
rect 140 256 141 257
rect 141 256 142 257
rect 142 256 143 257
rect 143 256 144 257
rect 144 256 145 257
rect 145 256 146 257
rect 146 256 147 257
rect 147 256 148 257
rect 148 256 149 257
rect 149 256 150 257
rect 150 256 151 257
rect 151 256 152 257
rect 152 256 153 257
rect 153 256 154 257
rect 154 256 155 257
rect 155 256 156 257
rect 156 256 157 257
rect 163 256 164 257
rect 164 256 165 257
rect 165 256 166 257
rect 166 256 167 257
rect 167 256 168 257
rect 168 256 169 257
rect 169 256 170 257
rect 170 256 171 257
rect 171 256 172 257
rect 172 256 173 257
rect 173 256 174 257
rect 174 256 175 257
rect 175 256 176 257
rect 176 256 177 257
rect 177 256 178 257
rect 178 256 179 257
rect 179 256 180 257
rect 180 256 181 257
rect 181 256 182 257
rect 182 256 183 257
rect 183 256 184 257
rect 184 256 185 257
rect 185 256 186 257
rect 186 256 187 257
rect 228 256 229 257
rect 229 256 230 257
rect 230 256 231 257
rect 231 256 232 257
rect 232 256 233 257
rect 233 256 234 257
rect 234 256 235 257
rect 235 256 236 257
rect 236 256 237 257
rect 237 256 238 257
rect 238 256 239 257
rect 239 256 240 257
rect 240 256 241 257
rect 241 256 242 257
rect 242 256 243 257
rect 243 256 244 257
rect 244 256 245 257
rect 245 256 246 257
rect 315 256 316 257
rect 316 256 317 257
rect 317 256 318 257
rect 348 256 349 257
rect 349 256 350 257
rect 350 256 351 257
rect 351 256 352 257
rect 352 256 353 257
rect 353 256 354 257
rect 354 256 355 257
rect 355 256 356 257
rect 356 256 357 257
rect 357 256 358 257
rect 383 256 384 257
rect 384 256 385 257
rect 385 256 386 257
rect 386 256 387 257
rect 387 256 388 257
rect 388 256 389 257
rect 389 256 390 257
rect 390 256 391 257
rect 63 255 64 256
rect 64 255 65 256
rect 65 255 66 256
rect 66 255 67 256
rect 67 255 68 256
rect 68 255 69 256
rect 69 255 70 256
rect 70 255 71 256
rect 71 255 72 256
rect 72 255 73 256
rect 73 255 74 256
rect 113 255 114 256
rect 114 255 115 256
rect 115 255 116 256
rect 116 255 117 256
rect 117 255 118 256
rect 118 255 119 256
rect 119 255 120 256
rect 120 255 121 256
rect 121 255 122 256
rect 122 255 123 256
rect 123 255 124 256
rect 124 255 125 256
rect 125 255 126 256
rect 126 255 127 256
rect 127 255 128 256
rect 128 255 129 256
rect 129 255 130 256
rect 130 255 131 256
rect 131 255 132 256
rect 132 255 133 256
rect 133 255 134 256
rect 134 255 135 256
rect 135 255 136 256
rect 136 255 137 256
rect 137 255 138 256
rect 138 255 139 256
rect 139 255 140 256
rect 140 255 141 256
rect 141 255 142 256
rect 142 255 143 256
rect 143 255 144 256
rect 144 255 145 256
rect 145 255 146 256
rect 146 255 147 256
rect 147 255 148 256
rect 148 255 149 256
rect 149 255 150 256
rect 150 255 151 256
rect 151 255 152 256
rect 152 255 153 256
rect 153 255 154 256
rect 158 255 159 256
rect 159 255 160 256
rect 160 255 161 256
rect 161 255 162 256
rect 162 255 163 256
rect 163 255 164 256
rect 164 255 165 256
rect 165 255 166 256
rect 166 255 167 256
rect 167 255 168 256
rect 168 255 169 256
rect 169 255 170 256
rect 170 255 171 256
rect 171 255 172 256
rect 172 255 173 256
rect 173 255 174 256
rect 174 255 175 256
rect 175 255 176 256
rect 176 255 177 256
rect 177 255 178 256
rect 178 255 179 256
rect 179 255 180 256
rect 180 255 181 256
rect 181 255 182 256
rect 182 255 183 256
rect 183 255 184 256
rect 184 255 185 256
rect 185 255 186 256
rect 186 255 187 256
rect 187 255 188 256
rect 227 255 228 256
rect 228 255 229 256
rect 229 255 230 256
rect 230 255 231 256
rect 231 255 232 256
rect 232 255 233 256
rect 233 255 234 256
rect 234 255 235 256
rect 235 255 236 256
rect 236 255 237 256
rect 237 255 238 256
rect 238 255 239 256
rect 239 255 240 256
rect 240 255 241 256
rect 241 255 242 256
rect 242 255 243 256
rect 243 255 244 256
rect 244 255 245 256
rect 245 255 246 256
rect 246 255 247 256
rect 247 255 248 256
rect 315 255 316 256
rect 316 255 317 256
rect 349 255 350 256
rect 350 255 351 256
rect 351 255 352 256
rect 352 255 353 256
rect 353 255 354 256
rect 354 255 355 256
rect 355 255 356 256
rect 356 255 357 256
rect 357 255 358 256
rect 383 255 384 256
rect 384 255 385 256
rect 385 255 386 256
rect 386 255 387 256
rect 387 255 388 256
rect 388 255 389 256
rect 389 255 390 256
rect 63 254 64 255
rect 64 254 65 255
rect 65 254 66 255
rect 66 254 67 255
rect 67 254 68 255
rect 68 254 69 255
rect 69 254 70 255
rect 70 254 71 255
rect 71 254 72 255
rect 72 254 73 255
rect 73 254 74 255
rect 113 254 114 255
rect 114 254 115 255
rect 115 254 116 255
rect 116 254 117 255
rect 117 254 118 255
rect 118 254 119 255
rect 119 254 120 255
rect 120 254 121 255
rect 121 254 122 255
rect 122 254 123 255
rect 123 254 124 255
rect 124 254 125 255
rect 125 254 126 255
rect 126 254 127 255
rect 127 254 128 255
rect 128 254 129 255
rect 129 254 130 255
rect 130 254 131 255
rect 131 254 132 255
rect 132 254 133 255
rect 133 254 134 255
rect 134 254 135 255
rect 135 254 136 255
rect 136 254 137 255
rect 137 254 138 255
rect 138 254 139 255
rect 139 254 140 255
rect 140 254 141 255
rect 141 254 142 255
rect 142 254 143 255
rect 143 254 144 255
rect 144 254 145 255
rect 145 254 146 255
rect 146 254 147 255
rect 147 254 148 255
rect 148 254 149 255
rect 149 254 150 255
rect 150 254 151 255
rect 151 254 152 255
rect 155 254 156 255
rect 156 254 157 255
rect 157 254 158 255
rect 158 254 159 255
rect 159 254 160 255
rect 160 254 161 255
rect 161 254 162 255
rect 162 254 163 255
rect 163 254 164 255
rect 164 254 165 255
rect 165 254 166 255
rect 166 254 167 255
rect 167 254 168 255
rect 168 254 169 255
rect 169 254 170 255
rect 170 254 171 255
rect 171 254 172 255
rect 172 254 173 255
rect 173 254 174 255
rect 174 254 175 255
rect 175 254 176 255
rect 176 254 177 255
rect 177 254 178 255
rect 178 254 179 255
rect 179 254 180 255
rect 180 254 181 255
rect 181 254 182 255
rect 182 254 183 255
rect 183 254 184 255
rect 184 254 185 255
rect 185 254 186 255
rect 186 254 187 255
rect 187 254 188 255
rect 227 254 228 255
rect 228 254 229 255
rect 229 254 230 255
rect 230 254 231 255
rect 231 254 232 255
rect 232 254 233 255
rect 233 254 234 255
rect 234 254 235 255
rect 235 254 236 255
rect 236 254 237 255
rect 237 254 238 255
rect 238 254 239 255
rect 239 254 240 255
rect 240 254 241 255
rect 241 254 242 255
rect 242 254 243 255
rect 243 254 244 255
rect 244 254 245 255
rect 245 254 246 255
rect 246 254 247 255
rect 247 254 248 255
rect 248 254 249 255
rect 249 254 250 255
rect 315 254 316 255
rect 316 254 317 255
rect 349 254 350 255
rect 350 254 351 255
rect 351 254 352 255
rect 352 254 353 255
rect 353 254 354 255
rect 354 254 355 255
rect 355 254 356 255
rect 356 254 357 255
rect 357 254 358 255
rect 382 254 383 255
rect 383 254 384 255
rect 384 254 385 255
rect 385 254 386 255
rect 386 254 387 255
rect 387 254 388 255
rect 388 254 389 255
rect 64 253 65 254
rect 65 253 66 254
rect 66 253 67 254
rect 67 253 68 254
rect 68 253 69 254
rect 69 253 70 254
rect 70 253 71 254
rect 71 253 72 254
rect 72 253 73 254
rect 73 253 74 254
rect 74 253 75 254
rect 114 253 115 254
rect 115 253 116 254
rect 116 253 117 254
rect 117 253 118 254
rect 118 253 119 254
rect 119 253 120 254
rect 120 253 121 254
rect 121 253 122 254
rect 122 253 123 254
rect 123 253 124 254
rect 124 253 125 254
rect 125 253 126 254
rect 126 253 127 254
rect 127 253 128 254
rect 128 253 129 254
rect 129 253 130 254
rect 130 253 131 254
rect 131 253 132 254
rect 132 253 133 254
rect 133 253 134 254
rect 134 253 135 254
rect 135 253 136 254
rect 136 253 137 254
rect 137 253 138 254
rect 138 253 139 254
rect 139 253 140 254
rect 140 253 141 254
rect 141 253 142 254
rect 142 253 143 254
rect 143 253 144 254
rect 144 253 145 254
rect 145 253 146 254
rect 146 253 147 254
rect 147 253 148 254
rect 148 253 149 254
rect 149 253 150 254
rect 152 253 153 254
rect 153 253 154 254
rect 154 253 155 254
rect 155 253 156 254
rect 156 253 157 254
rect 157 253 158 254
rect 158 253 159 254
rect 159 253 160 254
rect 160 253 161 254
rect 161 253 162 254
rect 162 253 163 254
rect 163 253 164 254
rect 164 253 165 254
rect 165 253 166 254
rect 166 253 167 254
rect 167 253 168 254
rect 168 253 169 254
rect 169 253 170 254
rect 170 253 171 254
rect 171 253 172 254
rect 172 253 173 254
rect 173 253 174 254
rect 174 253 175 254
rect 175 253 176 254
rect 176 253 177 254
rect 177 253 178 254
rect 178 253 179 254
rect 179 253 180 254
rect 180 253 181 254
rect 181 253 182 254
rect 182 253 183 254
rect 183 253 184 254
rect 184 253 185 254
rect 185 253 186 254
rect 186 253 187 254
rect 187 253 188 254
rect 226 253 227 254
rect 227 253 228 254
rect 228 253 229 254
rect 229 253 230 254
rect 230 253 231 254
rect 231 253 232 254
rect 232 253 233 254
rect 233 253 234 254
rect 234 253 235 254
rect 235 253 236 254
rect 236 253 237 254
rect 237 253 238 254
rect 238 253 239 254
rect 239 253 240 254
rect 240 253 241 254
rect 241 253 242 254
rect 242 253 243 254
rect 243 253 244 254
rect 244 253 245 254
rect 245 253 246 254
rect 246 253 247 254
rect 247 253 248 254
rect 248 253 249 254
rect 249 253 250 254
rect 250 253 251 254
rect 315 253 316 254
rect 316 253 317 254
rect 349 253 350 254
rect 350 253 351 254
rect 351 253 352 254
rect 352 253 353 254
rect 353 253 354 254
rect 354 253 355 254
rect 355 253 356 254
rect 356 253 357 254
rect 357 253 358 254
rect 381 253 382 254
rect 382 253 383 254
rect 383 253 384 254
rect 384 253 385 254
rect 385 253 386 254
rect 386 253 387 254
rect 387 253 388 254
rect 388 253 389 254
rect 65 252 66 253
rect 66 252 67 253
rect 67 252 68 253
rect 68 252 69 253
rect 69 252 70 253
rect 70 252 71 253
rect 71 252 72 253
rect 72 252 73 253
rect 73 252 74 253
rect 74 252 75 253
rect 75 252 76 253
rect 115 252 116 253
rect 116 252 117 253
rect 117 252 118 253
rect 118 252 119 253
rect 119 252 120 253
rect 120 252 121 253
rect 121 252 122 253
rect 122 252 123 253
rect 123 252 124 253
rect 124 252 125 253
rect 125 252 126 253
rect 126 252 127 253
rect 127 252 128 253
rect 128 252 129 253
rect 129 252 130 253
rect 130 252 131 253
rect 131 252 132 253
rect 132 252 133 253
rect 133 252 134 253
rect 134 252 135 253
rect 135 252 136 253
rect 136 252 137 253
rect 137 252 138 253
rect 138 252 139 253
rect 139 252 140 253
rect 140 252 141 253
rect 141 252 142 253
rect 142 252 143 253
rect 143 252 144 253
rect 144 252 145 253
rect 145 252 146 253
rect 146 252 147 253
rect 147 252 148 253
rect 150 252 151 253
rect 151 252 152 253
rect 152 252 153 253
rect 153 252 154 253
rect 154 252 155 253
rect 155 252 156 253
rect 156 252 157 253
rect 157 252 158 253
rect 158 252 159 253
rect 159 252 160 253
rect 160 252 161 253
rect 161 252 162 253
rect 162 252 163 253
rect 163 252 164 253
rect 164 252 165 253
rect 165 252 166 253
rect 166 252 167 253
rect 167 252 168 253
rect 168 252 169 253
rect 169 252 170 253
rect 170 252 171 253
rect 171 252 172 253
rect 172 252 173 253
rect 173 252 174 253
rect 174 252 175 253
rect 175 252 176 253
rect 176 252 177 253
rect 177 252 178 253
rect 178 252 179 253
rect 179 252 180 253
rect 180 252 181 253
rect 181 252 182 253
rect 182 252 183 253
rect 183 252 184 253
rect 184 252 185 253
rect 185 252 186 253
rect 186 252 187 253
rect 187 252 188 253
rect 225 252 226 253
rect 226 252 227 253
rect 227 252 228 253
rect 228 252 229 253
rect 229 252 230 253
rect 230 252 231 253
rect 231 252 232 253
rect 242 252 243 253
rect 243 252 244 253
rect 244 252 245 253
rect 245 252 246 253
rect 246 252 247 253
rect 247 252 248 253
rect 248 252 249 253
rect 249 252 250 253
rect 250 252 251 253
rect 251 252 252 253
rect 252 252 253 253
rect 315 252 316 253
rect 316 252 317 253
rect 350 252 351 253
rect 351 252 352 253
rect 352 252 353 253
rect 353 252 354 253
rect 354 252 355 253
rect 355 252 356 253
rect 356 252 357 253
rect 357 252 358 253
rect 358 252 359 253
rect 381 252 382 253
rect 382 252 383 253
rect 383 252 384 253
rect 384 252 385 253
rect 385 252 386 253
rect 386 252 387 253
rect 387 252 388 253
rect 65 251 66 252
rect 66 251 67 252
rect 67 251 68 252
rect 68 251 69 252
rect 69 251 70 252
rect 70 251 71 252
rect 71 251 72 252
rect 72 251 73 252
rect 73 251 74 252
rect 74 251 75 252
rect 75 251 76 252
rect 76 251 77 252
rect 115 251 116 252
rect 116 251 117 252
rect 117 251 118 252
rect 118 251 119 252
rect 119 251 120 252
rect 120 251 121 252
rect 121 251 122 252
rect 122 251 123 252
rect 123 251 124 252
rect 124 251 125 252
rect 125 251 126 252
rect 126 251 127 252
rect 127 251 128 252
rect 128 251 129 252
rect 129 251 130 252
rect 130 251 131 252
rect 131 251 132 252
rect 132 251 133 252
rect 133 251 134 252
rect 134 251 135 252
rect 135 251 136 252
rect 136 251 137 252
rect 137 251 138 252
rect 138 251 139 252
rect 139 251 140 252
rect 140 251 141 252
rect 141 251 142 252
rect 142 251 143 252
rect 143 251 144 252
rect 144 251 145 252
rect 145 251 146 252
rect 146 251 147 252
rect 147 251 148 252
rect 148 251 149 252
rect 149 251 150 252
rect 150 251 151 252
rect 151 251 152 252
rect 152 251 153 252
rect 153 251 154 252
rect 154 251 155 252
rect 155 251 156 252
rect 156 251 157 252
rect 157 251 158 252
rect 158 251 159 252
rect 159 251 160 252
rect 160 251 161 252
rect 161 251 162 252
rect 162 251 163 252
rect 163 251 164 252
rect 164 251 165 252
rect 165 251 166 252
rect 166 251 167 252
rect 167 251 168 252
rect 168 251 169 252
rect 169 251 170 252
rect 170 251 171 252
rect 171 251 172 252
rect 172 251 173 252
rect 173 251 174 252
rect 174 251 175 252
rect 175 251 176 252
rect 176 251 177 252
rect 177 251 178 252
rect 178 251 179 252
rect 179 251 180 252
rect 180 251 181 252
rect 181 251 182 252
rect 182 251 183 252
rect 183 251 184 252
rect 184 251 185 252
rect 185 251 186 252
rect 186 251 187 252
rect 187 251 188 252
rect 223 251 224 252
rect 224 251 225 252
rect 225 251 226 252
rect 226 251 227 252
rect 227 251 228 252
rect 228 251 229 252
rect 229 251 230 252
rect 230 251 231 252
rect 231 251 232 252
rect 232 251 233 252
rect 233 251 234 252
rect 234 251 235 252
rect 235 251 236 252
rect 236 251 237 252
rect 237 251 238 252
rect 244 251 245 252
rect 245 251 246 252
rect 246 251 247 252
rect 247 251 248 252
rect 248 251 249 252
rect 249 251 250 252
rect 250 251 251 252
rect 251 251 252 252
rect 252 251 253 252
rect 253 251 254 252
rect 314 251 315 252
rect 315 251 316 252
rect 316 251 317 252
rect 350 251 351 252
rect 351 251 352 252
rect 352 251 353 252
rect 353 251 354 252
rect 354 251 355 252
rect 355 251 356 252
rect 356 251 357 252
rect 357 251 358 252
rect 358 251 359 252
rect 380 251 381 252
rect 381 251 382 252
rect 382 251 383 252
rect 383 251 384 252
rect 384 251 385 252
rect 385 251 386 252
rect 386 251 387 252
rect 387 251 388 252
rect 66 250 67 251
rect 67 250 68 251
rect 68 250 69 251
rect 69 250 70 251
rect 70 250 71 251
rect 71 250 72 251
rect 72 250 73 251
rect 73 250 74 251
rect 74 250 75 251
rect 75 250 76 251
rect 76 250 77 251
rect 77 250 78 251
rect 116 250 117 251
rect 117 250 118 251
rect 118 250 119 251
rect 119 250 120 251
rect 120 250 121 251
rect 121 250 122 251
rect 122 250 123 251
rect 123 250 124 251
rect 124 250 125 251
rect 125 250 126 251
rect 126 250 127 251
rect 127 250 128 251
rect 128 250 129 251
rect 129 250 130 251
rect 130 250 131 251
rect 131 250 132 251
rect 132 250 133 251
rect 133 250 134 251
rect 134 250 135 251
rect 135 250 136 251
rect 136 250 137 251
rect 137 250 138 251
rect 138 250 139 251
rect 139 250 140 251
rect 140 250 141 251
rect 141 250 142 251
rect 142 250 143 251
rect 143 250 144 251
rect 144 250 145 251
rect 145 250 146 251
rect 146 250 147 251
rect 147 250 148 251
rect 148 250 149 251
rect 149 250 150 251
rect 150 250 151 251
rect 151 250 152 251
rect 152 250 153 251
rect 153 250 154 251
rect 154 250 155 251
rect 155 250 156 251
rect 156 250 157 251
rect 157 250 158 251
rect 158 250 159 251
rect 159 250 160 251
rect 160 250 161 251
rect 161 250 162 251
rect 162 250 163 251
rect 163 250 164 251
rect 164 250 165 251
rect 165 250 166 251
rect 166 250 167 251
rect 167 250 168 251
rect 168 250 169 251
rect 169 250 170 251
rect 170 250 171 251
rect 171 250 172 251
rect 172 250 173 251
rect 173 250 174 251
rect 174 250 175 251
rect 175 250 176 251
rect 176 250 177 251
rect 177 250 178 251
rect 178 250 179 251
rect 179 250 180 251
rect 180 250 181 251
rect 181 250 182 251
rect 182 250 183 251
rect 183 250 184 251
rect 184 250 185 251
rect 185 250 186 251
rect 186 250 187 251
rect 187 250 188 251
rect 220 250 221 251
rect 221 250 222 251
rect 222 250 223 251
rect 223 250 224 251
rect 224 250 225 251
rect 225 250 226 251
rect 226 250 227 251
rect 227 250 228 251
rect 228 250 229 251
rect 229 250 230 251
rect 230 250 231 251
rect 231 250 232 251
rect 232 250 233 251
rect 233 250 234 251
rect 234 250 235 251
rect 235 250 236 251
rect 236 250 237 251
rect 237 250 238 251
rect 238 250 239 251
rect 239 250 240 251
rect 240 250 241 251
rect 241 250 242 251
rect 247 250 248 251
rect 248 250 249 251
rect 249 250 250 251
rect 250 250 251 251
rect 251 250 252 251
rect 252 250 253 251
rect 253 250 254 251
rect 254 250 255 251
rect 314 250 315 251
rect 315 250 316 251
rect 316 250 317 251
rect 350 250 351 251
rect 351 250 352 251
rect 352 250 353 251
rect 353 250 354 251
rect 354 250 355 251
rect 355 250 356 251
rect 356 250 357 251
rect 357 250 358 251
rect 358 250 359 251
rect 359 250 360 251
rect 379 250 380 251
rect 380 250 381 251
rect 381 250 382 251
rect 382 250 383 251
rect 383 250 384 251
rect 384 250 385 251
rect 385 250 386 251
rect 386 250 387 251
rect 67 249 68 250
rect 68 249 69 250
rect 69 249 70 250
rect 70 249 71 250
rect 71 249 72 250
rect 72 249 73 250
rect 73 249 74 250
rect 74 249 75 250
rect 75 249 76 250
rect 76 249 77 250
rect 77 249 78 250
rect 78 249 79 250
rect 117 249 118 250
rect 118 249 119 250
rect 119 249 120 250
rect 120 249 121 250
rect 121 249 122 250
rect 122 249 123 250
rect 123 249 124 250
rect 124 249 125 250
rect 125 249 126 250
rect 126 249 127 250
rect 127 249 128 250
rect 128 249 129 250
rect 129 249 130 250
rect 130 249 131 250
rect 131 249 132 250
rect 132 249 133 250
rect 133 249 134 250
rect 134 249 135 250
rect 135 249 136 250
rect 136 249 137 250
rect 137 249 138 250
rect 138 249 139 250
rect 139 249 140 250
rect 140 249 141 250
rect 141 249 142 250
rect 142 249 143 250
rect 143 249 144 250
rect 144 249 145 250
rect 145 249 146 250
rect 146 249 147 250
rect 147 249 148 250
rect 148 249 149 250
rect 149 249 150 250
rect 150 249 151 250
rect 151 249 152 250
rect 152 249 153 250
rect 153 249 154 250
rect 154 249 155 250
rect 155 249 156 250
rect 156 249 157 250
rect 157 249 158 250
rect 158 249 159 250
rect 159 249 160 250
rect 160 249 161 250
rect 161 249 162 250
rect 162 249 163 250
rect 163 249 164 250
rect 164 249 165 250
rect 165 249 166 250
rect 166 249 167 250
rect 167 249 168 250
rect 168 249 169 250
rect 169 249 170 250
rect 170 249 171 250
rect 171 249 172 250
rect 172 249 173 250
rect 173 249 174 250
rect 174 249 175 250
rect 175 249 176 250
rect 176 249 177 250
rect 177 249 178 250
rect 178 249 179 250
rect 179 249 180 250
rect 180 249 181 250
rect 181 249 182 250
rect 182 249 183 250
rect 183 249 184 250
rect 184 249 185 250
rect 185 249 186 250
rect 186 249 187 250
rect 187 249 188 250
rect 216 249 217 250
rect 217 249 218 250
rect 218 249 219 250
rect 219 249 220 250
rect 220 249 221 250
rect 221 249 222 250
rect 222 249 223 250
rect 223 249 224 250
rect 224 249 225 250
rect 225 249 226 250
rect 226 249 227 250
rect 233 249 234 250
rect 234 249 235 250
rect 235 249 236 250
rect 236 249 237 250
rect 237 249 238 250
rect 238 249 239 250
rect 239 249 240 250
rect 240 249 241 250
rect 241 249 242 250
rect 242 249 243 250
rect 243 249 244 250
rect 248 249 249 250
rect 249 249 250 250
rect 250 249 251 250
rect 251 249 252 250
rect 252 249 253 250
rect 253 249 254 250
rect 254 249 255 250
rect 255 249 256 250
rect 256 249 257 250
rect 314 249 315 250
rect 315 249 316 250
rect 316 249 317 250
rect 350 249 351 250
rect 351 249 352 250
rect 352 249 353 250
rect 353 249 354 250
rect 354 249 355 250
rect 355 249 356 250
rect 356 249 357 250
rect 357 249 358 250
rect 358 249 359 250
rect 359 249 360 250
rect 360 249 361 250
rect 378 249 379 250
rect 379 249 380 250
rect 380 249 381 250
rect 381 249 382 250
rect 382 249 383 250
rect 383 249 384 250
rect 384 249 385 250
rect 385 249 386 250
rect 68 248 69 249
rect 69 248 70 249
rect 70 248 71 249
rect 71 248 72 249
rect 72 248 73 249
rect 73 248 74 249
rect 74 248 75 249
rect 75 248 76 249
rect 76 248 77 249
rect 77 248 78 249
rect 78 248 79 249
rect 79 248 80 249
rect 118 248 119 249
rect 119 248 120 249
rect 120 248 121 249
rect 121 248 122 249
rect 122 248 123 249
rect 123 248 124 249
rect 124 248 125 249
rect 125 248 126 249
rect 126 248 127 249
rect 127 248 128 249
rect 128 248 129 249
rect 129 248 130 249
rect 130 248 131 249
rect 131 248 132 249
rect 132 248 133 249
rect 133 248 134 249
rect 134 248 135 249
rect 135 248 136 249
rect 136 248 137 249
rect 137 248 138 249
rect 138 248 139 249
rect 139 248 140 249
rect 140 248 141 249
rect 141 248 142 249
rect 142 248 143 249
rect 143 248 144 249
rect 144 248 145 249
rect 145 248 146 249
rect 146 248 147 249
rect 147 248 148 249
rect 148 248 149 249
rect 149 248 150 249
rect 150 248 151 249
rect 151 248 152 249
rect 152 248 153 249
rect 153 248 154 249
rect 154 248 155 249
rect 155 248 156 249
rect 156 248 157 249
rect 157 248 158 249
rect 158 248 159 249
rect 159 248 160 249
rect 160 248 161 249
rect 161 248 162 249
rect 162 248 163 249
rect 163 248 164 249
rect 164 248 165 249
rect 165 248 166 249
rect 166 248 167 249
rect 167 248 168 249
rect 168 248 169 249
rect 169 248 170 249
rect 170 248 171 249
rect 171 248 172 249
rect 172 248 173 249
rect 173 248 174 249
rect 174 248 175 249
rect 175 248 176 249
rect 176 248 177 249
rect 177 248 178 249
rect 178 248 179 249
rect 179 248 180 249
rect 180 248 181 249
rect 181 248 182 249
rect 182 248 183 249
rect 183 248 184 249
rect 184 248 185 249
rect 185 248 186 249
rect 186 248 187 249
rect 187 248 188 249
rect 215 248 216 249
rect 216 248 217 249
rect 217 248 218 249
rect 218 248 219 249
rect 219 248 220 249
rect 220 248 221 249
rect 221 248 222 249
rect 222 248 223 249
rect 223 248 224 249
rect 224 248 225 249
rect 226 248 227 249
rect 227 248 228 249
rect 236 248 237 249
rect 237 248 238 249
rect 238 248 239 249
rect 239 248 240 249
rect 240 248 241 249
rect 241 248 242 249
rect 242 248 243 249
rect 243 248 244 249
rect 244 248 245 249
rect 245 248 246 249
rect 250 248 251 249
rect 251 248 252 249
rect 252 248 253 249
rect 253 248 254 249
rect 254 248 255 249
rect 255 248 256 249
rect 256 248 257 249
rect 257 248 258 249
rect 292 248 293 249
rect 314 248 315 249
rect 315 248 316 249
rect 316 248 317 249
rect 350 248 351 249
rect 351 248 352 249
rect 352 248 353 249
rect 353 248 354 249
rect 354 248 355 249
rect 355 248 356 249
rect 356 248 357 249
rect 357 248 358 249
rect 358 248 359 249
rect 359 248 360 249
rect 360 248 361 249
rect 378 248 379 249
rect 379 248 380 249
rect 380 248 381 249
rect 381 248 382 249
rect 382 248 383 249
rect 383 248 384 249
rect 384 248 385 249
rect 385 248 386 249
rect 69 247 70 248
rect 70 247 71 248
rect 71 247 72 248
rect 72 247 73 248
rect 73 247 74 248
rect 74 247 75 248
rect 75 247 76 248
rect 76 247 77 248
rect 77 247 78 248
rect 78 247 79 248
rect 79 247 80 248
rect 80 247 81 248
rect 120 247 121 248
rect 121 247 122 248
rect 122 247 123 248
rect 123 247 124 248
rect 124 247 125 248
rect 125 247 126 248
rect 126 247 127 248
rect 127 247 128 248
rect 128 247 129 248
rect 129 247 130 248
rect 130 247 131 248
rect 131 247 132 248
rect 132 247 133 248
rect 133 247 134 248
rect 134 247 135 248
rect 135 247 136 248
rect 136 247 137 248
rect 137 247 138 248
rect 138 247 139 248
rect 139 247 140 248
rect 140 247 141 248
rect 141 247 142 248
rect 142 247 143 248
rect 143 247 144 248
rect 144 247 145 248
rect 145 247 146 248
rect 146 247 147 248
rect 147 247 148 248
rect 148 247 149 248
rect 149 247 150 248
rect 150 247 151 248
rect 151 247 152 248
rect 152 247 153 248
rect 153 247 154 248
rect 154 247 155 248
rect 155 247 156 248
rect 156 247 157 248
rect 157 247 158 248
rect 158 247 159 248
rect 159 247 160 248
rect 160 247 161 248
rect 161 247 162 248
rect 162 247 163 248
rect 163 247 164 248
rect 164 247 165 248
rect 165 247 166 248
rect 166 247 167 248
rect 167 247 168 248
rect 168 247 169 248
rect 169 247 170 248
rect 170 247 171 248
rect 171 247 172 248
rect 172 247 173 248
rect 173 247 174 248
rect 174 247 175 248
rect 175 247 176 248
rect 176 247 177 248
rect 177 247 178 248
rect 178 247 179 248
rect 179 247 180 248
rect 180 247 181 248
rect 181 247 182 248
rect 182 247 183 248
rect 183 247 184 248
rect 184 247 185 248
rect 185 247 186 248
rect 186 247 187 248
rect 187 247 188 248
rect 215 247 216 248
rect 216 247 217 248
rect 217 247 218 248
rect 218 247 219 248
rect 219 247 220 248
rect 220 247 221 248
rect 221 247 222 248
rect 222 247 223 248
rect 223 247 224 248
rect 224 247 225 248
rect 225 247 226 248
rect 226 247 227 248
rect 227 247 228 248
rect 228 247 229 248
rect 229 247 230 248
rect 230 247 231 248
rect 231 247 232 248
rect 232 247 233 248
rect 239 247 240 248
rect 240 247 241 248
rect 241 247 242 248
rect 242 247 243 248
rect 243 247 244 248
rect 244 247 245 248
rect 245 247 246 248
rect 246 247 247 248
rect 247 247 248 248
rect 251 247 252 248
rect 252 247 253 248
rect 253 247 254 248
rect 254 247 255 248
rect 255 247 256 248
rect 256 247 257 248
rect 257 247 258 248
rect 258 247 259 248
rect 290 247 291 248
rect 291 247 292 248
rect 292 247 293 248
rect 314 247 315 248
rect 315 247 316 248
rect 316 247 317 248
rect 350 247 351 248
rect 351 247 352 248
rect 352 247 353 248
rect 356 247 357 248
rect 357 247 358 248
rect 358 247 359 248
rect 359 247 360 248
rect 360 247 361 248
rect 361 247 362 248
rect 377 247 378 248
rect 378 247 379 248
rect 379 247 380 248
rect 380 247 381 248
rect 381 247 382 248
rect 382 247 383 248
rect 383 247 384 248
rect 384 247 385 248
rect 385 247 386 248
rect 69 246 70 247
rect 70 246 71 247
rect 71 246 72 247
rect 72 246 73 247
rect 73 246 74 247
rect 74 246 75 247
rect 75 246 76 247
rect 76 246 77 247
rect 77 246 78 247
rect 78 246 79 247
rect 79 246 80 247
rect 80 246 81 247
rect 81 246 82 247
rect 121 246 122 247
rect 122 246 123 247
rect 123 246 124 247
rect 124 246 125 247
rect 125 246 126 247
rect 126 246 127 247
rect 127 246 128 247
rect 128 246 129 247
rect 129 246 130 247
rect 130 246 131 247
rect 131 246 132 247
rect 132 246 133 247
rect 133 246 134 247
rect 134 246 135 247
rect 135 246 136 247
rect 136 246 137 247
rect 137 246 138 247
rect 138 246 139 247
rect 139 246 140 247
rect 140 246 141 247
rect 141 246 142 247
rect 142 246 143 247
rect 143 246 144 247
rect 144 246 145 247
rect 145 246 146 247
rect 146 246 147 247
rect 147 246 148 247
rect 148 246 149 247
rect 149 246 150 247
rect 150 246 151 247
rect 151 246 152 247
rect 152 246 153 247
rect 153 246 154 247
rect 154 246 155 247
rect 155 246 156 247
rect 156 246 157 247
rect 157 246 158 247
rect 158 246 159 247
rect 159 246 160 247
rect 160 246 161 247
rect 161 246 162 247
rect 162 246 163 247
rect 163 246 164 247
rect 164 246 165 247
rect 165 246 166 247
rect 166 246 167 247
rect 167 246 168 247
rect 168 246 169 247
rect 169 246 170 247
rect 170 246 171 247
rect 171 246 172 247
rect 172 246 173 247
rect 173 246 174 247
rect 174 246 175 247
rect 175 246 176 247
rect 176 246 177 247
rect 177 246 178 247
rect 178 246 179 247
rect 179 246 180 247
rect 180 246 181 247
rect 181 246 182 247
rect 182 246 183 247
rect 183 246 184 247
rect 184 246 185 247
rect 185 246 186 247
rect 186 246 187 247
rect 187 246 188 247
rect 215 246 216 247
rect 216 246 217 247
rect 217 246 218 247
rect 218 246 219 247
rect 219 246 220 247
rect 220 246 221 247
rect 221 246 222 247
rect 222 246 223 247
rect 223 246 224 247
rect 224 246 225 247
rect 225 246 226 247
rect 226 246 227 247
rect 227 246 228 247
rect 228 246 229 247
rect 229 246 230 247
rect 230 246 231 247
rect 231 246 232 247
rect 232 246 233 247
rect 233 246 234 247
rect 234 246 235 247
rect 235 246 236 247
rect 241 246 242 247
rect 242 246 243 247
rect 243 246 244 247
rect 244 246 245 247
rect 245 246 246 247
rect 246 246 247 247
rect 247 246 248 247
rect 248 246 249 247
rect 249 246 250 247
rect 253 246 254 247
rect 254 246 255 247
rect 255 246 256 247
rect 256 246 257 247
rect 257 246 258 247
rect 258 246 259 247
rect 259 246 260 247
rect 260 246 261 247
rect 288 246 289 247
rect 289 246 290 247
rect 290 246 291 247
rect 291 246 292 247
rect 314 246 315 247
rect 315 246 316 247
rect 316 246 317 247
rect 350 246 351 247
rect 351 246 352 247
rect 358 246 359 247
rect 359 246 360 247
rect 360 246 361 247
rect 361 246 362 247
rect 376 246 377 247
rect 377 246 378 247
rect 378 246 379 247
rect 379 246 380 247
rect 380 246 381 247
rect 381 246 382 247
rect 382 246 383 247
rect 383 246 384 247
rect 384 246 385 247
rect 385 246 386 247
rect 386 246 387 247
rect 387 246 388 247
rect 70 245 71 246
rect 71 245 72 246
rect 72 245 73 246
rect 73 245 74 246
rect 74 245 75 246
rect 75 245 76 246
rect 76 245 77 246
rect 77 245 78 246
rect 78 245 79 246
rect 79 245 80 246
rect 80 245 81 246
rect 81 245 82 246
rect 82 245 83 246
rect 124 245 125 246
rect 125 245 126 246
rect 126 245 127 246
rect 127 245 128 246
rect 128 245 129 246
rect 129 245 130 246
rect 130 245 131 246
rect 131 245 132 246
rect 132 245 133 246
rect 133 245 134 246
rect 134 245 135 246
rect 135 245 136 246
rect 136 245 137 246
rect 137 245 138 246
rect 138 245 139 246
rect 139 245 140 246
rect 140 245 141 246
rect 141 245 142 246
rect 142 245 143 246
rect 143 245 144 246
rect 144 245 145 246
rect 145 245 146 246
rect 146 245 147 246
rect 147 245 148 246
rect 148 245 149 246
rect 149 245 150 246
rect 150 245 151 246
rect 151 245 152 246
rect 152 245 153 246
rect 153 245 154 246
rect 154 245 155 246
rect 155 245 156 246
rect 156 245 157 246
rect 157 245 158 246
rect 158 245 159 246
rect 159 245 160 246
rect 160 245 161 246
rect 161 245 162 246
rect 162 245 163 246
rect 163 245 164 246
rect 164 245 165 246
rect 165 245 166 246
rect 166 245 167 246
rect 167 245 168 246
rect 168 245 169 246
rect 169 245 170 246
rect 170 245 171 246
rect 171 245 172 246
rect 172 245 173 246
rect 173 245 174 246
rect 174 245 175 246
rect 175 245 176 246
rect 176 245 177 246
rect 177 245 178 246
rect 178 245 179 246
rect 179 245 180 246
rect 180 245 181 246
rect 181 245 182 246
rect 182 245 183 246
rect 183 245 184 246
rect 184 245 185 246
rect 185 245 186 246
rect 186 245 187 246
rect 187 245 188 246
rect 215 245 216 246
rect 216 245 217 246
rect 217 245 218 246
rect 218 245 219 246
rect 219 245 220 246
rect 220 245 221 246
rect 221 245 222 246
rect 222 245 223 246
rect 223 245 224 246
rect 224 245 225 246
rect 225 245 226 246
rect 226 245 227 246
rect 227 245 228 246
rect 228 245 229 246
rect 229 245 230 246
rect 230 245 231 246
rect 231 245 232 246
rect 232 245 233 246
rect 233 245 234 246
rect 234 245 235 246
rect 235 245 236 246
rect 236 245 237 246
rect 237 245 238 246
rect 242 245 243 246
rect 243 245 244 246
rect 244 245 245 246
rect 245 245 246 246
rect 246 245 247 246
rect 247 245 248 246
rect 248 245 249 246
rect 249 245 250 246
rect 250 245 251 246
rect 251 245 252 246
rect 254 245 255 246
rect 255 245 256 246
rect 256 245 257 246
rect 257 245 258 246
rect 258 245 259 246
rect 259 245 260 246
rect 260 245 261 246
rect 261 245 262 246
rect 262 245 263 246
rect 286 245 287 246
rect 287 245 288 246
rect 288 245 289 246
rect 289 245 290 246
rect 290 245 291 246
rect 314 245 315 246
rect 315 245 316 246
rect 316 245 317 246
rect 317 245 318 246
rect 350 245 351 246
rect 351 245 352 246
rect 360 245 361 246
rect 361 245 362 246
rect 362 245 363 246
rect 375 245 376 246
rect 376 245 377 246
rect 377 245 378 246
rect 378 245 379 246
rect 379 245 380 246
rect 380 245 381 246
rect 381 245 382 246
rect 382 245 383 246
rect 383 245 384 246
rect 384 245 385 246
rect 385 245 386 246
rect 386 245 387 246
rect 387 245 388 246
rect 388 245 389 246
rect 389 245 390 246
rect 71 244 72 245
rect 72 244 73 245
rect 73 244 74 245
rect 74 244 75 245
rect 75 244 76 245
rect 76 244 77 245
rect 77 244 78 245
rect 78 244 79 245
rect 79 244 80 245
rect 80 244 81 245
rect 81 244 82 245
rect 82 244 83 245
rect 83 244 84 245
rect 123 244 124 245
rect 124 244 125 245
rect 125 244 126 245
rect 126 244 127 245
rect 127 244 128 245
rect 128 244 129 245
rect 129 244 130 245
rect 130 244 131 245
rect 131 244 132 245
rect 132 244 133 245
rect 133 244 134 245
rect 134 244 135 245
rect 135 244 136 245
rect 136 244 137 245
rect 137 244 138 245
rect 138 244 139 245
rect 139 244 140 245
rect 140 244 141 245
rect 141 244 142 245
rect 142 244 143 245
rect 143 244 144 245
rect 144 244 145 245
rect 145 244 146 245
rect 146 244 147 245
rect 147 244 148 245
rect 148 244 149 245
rect 149 244 150 245
rect 150 244 151 245
rect 151 244 152 245
rect 152 244 153 245
rect 153 244 154 245
rect 154 244 155 245
rect 155 244 156 245
rect 156 244 157 245
rect 157 244 158 245
rect 158 244 159 245
rect 159 244 160 245
rect 160 244 161 245
rect 161 244 162 245
rect 162 244 163 245
rect 163 244 164 245
rect 164 244 165 245
rect 165 244 166 245
rect 166 244 167 245
rect 167 244 168 245
rect 168 244 169 245
rect 169 244 170 245
rect 170 244 171 245
rect 171 244 172 245
rect 172 244 173 245
rect 173 244 174 245
rect 174 244 175 245
rect 175 244 176 245
rect 176 244 177 245
rect 177 244 178 245
rect 178 244 179 245
rect 179 244 180 245
rect 180 244 181 245
rect 181 244 182 245
rect 182 244 183 245
rect 183 244 184 245
rect 184 244 185 245
rect 185 244 186 245
rect 186 244 187 245
rect 187 244 188 245
rect 214 244 215 245
rect 215 244 216 245
rect 216 244 217 245
rect 217 244 218 245
rect 218 244 219 245
rect 219 244 220 245
rect 220 244 221 245
rect 221 244 222 245
rect 222 244 223 245
rect 223 244 224 245
rect 224 244 225 245
rect 225 244 226 245
rect 226 244 227 245
rect 227 244 228 245
rect 228 244 229 245
rect 229 244 230 245
rect 230 244 231 245
rect 231 244 232 245
rect 232 244 233 245
rect 233 244 234 245
rect 234 244 235 245
rect 235 244 236 245
rect 236 244 237 245
rect 237 244 238 245
rect 238 244 239 245
rect 239 244 240 245
rect 244 244 245 245
rect 245 244 246 245
rect 246 244 247 245
rect 247 244 248 245
rect 248 244 249 245
rect 249 244 250 245
rect 250 244 251 245
rect 251 244 252 245
rect 252 244 253 245
rect 255 244 256 245
rect 256 244 257 245
rect 257 244 258 245
rect 258 244 259 245
rect 259 244 260 245
rect 260 244 261 245
rect 261 244 262 245
rect 262 244 263 245
rect 263 244 264 245
rect 264 244 265 245
rect 283 244 284 245
rect 284 244 285 245
rect 285 244 286 245
rect 286 244 287 245
rect 287 244 288 245
rect 288 244 289 245
rect 289 244 290 245
rect 290 244 291 245
rect 314 244 315 245
rect 315 244 316 245
rect 316 244 317 245
rect 317 244 318 245
rect 350 244 351 245
rect 361 244 362 245
rect 362 244 363 245
rect 374 244 375 245
rect 375 244 376 245
rect 376 244 377 245
rect 377 244 378 245
rect 378 244 379 245
rect 379 244 380 245
rect 380 244 381 245
rect 381 244 382 245
rect 382 244 383 245
rect 383 244 384 245
rect 384 244 385 245
rect 385 244 386 245
rect 386 244 387 245
rect 387 244 388 245
rect 388 244 389 245
rect 389 244 390 245
rect 390 244 391 245
rect 391 244 392 245
rect 392 244 393 245
rect 72 243 73 244
rect 73 243 74 244
rect 74 243 75 244
rect 75 243 76 244
rect 76 243 77 244
rect 77 243 78 244
rect 78 243 79 244
rect 79 243 80 244
rect 80 243 81 244
rect 81 243 82 244
rect 82 243 83 244
rect 83 243 84 244
rect 84 243 85 244
rect 85 243 86 244
rect 120 243 121 244
rect 121 243 122 244
rect 122 243 123 244
rect 123 243 124 244
rect 124 243 125 244
rect 125 243 126 244
rect 126 243 127 244
rect 127 243 128 244
rect 128 243 129 244
rect 129 243 130 244
rect 130 243 131 244
rect 131 243 132 244
rect 132 243 133 244
rect 133 243 134 244
rect 134 243 135 244
rect 135 243 136 244
rect 136 243 137 244
rect 137 243 138 244
rect 138 243 139 244
rect 139 243 140 244
rect 140 243 141 244
rect 141 243 142 244
rect 142 243 143 244
rect 143 243 144 244
rect 144 243 145 244
rect 145 243 146 244
rect 146 243 147 244
rect 147 243 148 244
rect 148 243 149 244
rect 149 243 150 244
rect 150 243 151 244
rect 151 243 152 244
rect 152 243 153 244
rect 153 243 154 244
rect 154 243 155 244
rect 155 243 156 244
rect 156 243 157 244
rect 157 243 158 244
rect 158 243 159 244
rect 159 243 160 244
rect 160 243 161 244
rect 161 243 162 244
rect 162 243 163 244
rect 163 243 164 244
rect 164 243 165 244
rect 165 243 166 244
rect 166 243 167 244
rect 167 243 168 244
rect 168 243 169 244
rect 169 243 170 244
rect 170 243 171 244
rect 171 243 172 244
rect 172 243 173 244
rect 173 243 174 244
rect 174 243 175 244
rect 175 243 176 244
rect 176 243 177 244
rect 177 243 178 244
rect 178 243 179 244
rect 179 243 180 244
rect 180 243 181 244
rect 181 243 182 244
rect 182 243 183 244
rect 183 243 184 244
rect 184 243 185 244
rect 185 243 186 244
rect 186 243 187 244
rect 187 243 188 244
rect 214 243 215 244
rect 215 243 216 244
rect 216 243 217 244
rect 217 243 218 244
rect 218 243 219 244
rect 219 243 220 244
rect 220 243 221 244
rect 221 243 222 244
rect 222 243 223 244
rect 223 243 224 244
rect 224 243 225 244
rect 225 243 226 244
rect 226 243 227 244
rect 227 243 228 244
rect 228 243 229 244
rect 229 243 230 244
rect 230 243 231 244
rect 231 243 232 244
rect 232 243 233 244
rect 233 243 234 244
rect 234 243 235 244
rect 235 243 236 244
rect 236 243 237 244
rect 237 243 238 244
rect 238 243 239 244
rect 239 243 240 244
rect 240 243 241 244
rect 241 243 242 244
rect 245 243 246 244
rect 246 243 247 244
rect 247 243 248 244
rect 248 243 249 244
rect 249 243 250 244
rect 250 243 251 244
rect 251 243 252 244
rect 252 243 253 244
rect 253 243 254 244
rect 254 243 255 244
rect 256 243 257 244
rect 257 243 258 244
rect 258 243 259 244
rect 259 243 260 244
rect 260 243 261 244
rect 261 243 262 244
rect 262 243 263 244
rect 263 243 264 244
rect 264 243 265 244
rect 265 243 266 244
rect 266 243 267 244
rect 267 243 268 244
rect 280 243 281 244
rect 281 243 282 244
rect 282 243 283 244
rect 283 243 284 244
rect 284 243 285 244
rect 285 243 286 244
rect 286 243 287 244
rect 287 243 288 244
rect 288 243 289 244
rect 289 243 290 244
rect 315 243 316 244
rect 316 243 317 244
rect 317 243 318 244
rect 318 243 319 244
rect 362 243 363 244
rect 373 243 374 244
rect 374 243 375 244
rect 375 243 376 244
rect 376 243 377 244
rect 377 243 378 244
rect 378 243 379 244
rect 379 243 380 244
rect 380 243 381 244
rect 381 243 382 244
rect 382 243 383 244
rect 383 243 384 244
rect 384 243 385 244
rect 385 243 386 244
rect 386 243 387 244
rect 387 243 388 244
rect 388 243 389 244
rect 389 243 390 244
rect 390 243 391 244
rect 391 243 392 244
rect 392 243 393 244
rect 393 243 394 244
rect 394 243 395 244
rect 395 243 396 244
rect 73 242 74 243
rect 74 242 75 243
rect 75 242 76 243
rect 76 242 77 243
rect 77 242 78 243
rect 78 242 79 243
rect 79 242 80 243
rect 80 242 81 243
rect 81 242 82 243
rect 82 242 83 243
rect 83 242 84 243
rect 84 242 85 243
rect 85 242 86 243
rect 86 242 87 243
rect 96 242 97 243
rect 97 242 98 243
rect 98 242 99 243
rect 118 242 119 243
rect 119 242 120 243
rect 120 242 121 243
rect 121 242 122 243
rect 122 242 123 243
rect 123 242 124 243
rect 124 242 125 243
rect 125 242 126 243
rect 126 242 127 243
rect 127 242 128 243
rect 128 242 129 243
rect 129 242 130 243
rect 130 242 131 243
rect 131 242 132 243
rect 132 242 133 243
rect 133 242 134 243
rect 134 242 135 243
rect 135 242 136 243
rect 136 242 137 243
rect 137 242 138 243
rect 138 242 139 243
rect 139 242 140 243
rect 140 242 141 243
rect 141 242 142 243
rect 142 242 143 243
rect 143 242 144 243
rect 144 242 145 243
rect 145 242 146 243
rect 146 242 147 243
rect 147 242 148 243
rect 148 242 149 243
rect 149 242 150 243
rect 150 242 151 243
rect 151 242 152 243
rect 152 242 153 243
rect 153 242 154 243
rect 154 242 155 243
rect 155 242 156 243
rect 156 242 157 243
rect 157 242 158 243
rect 158 242 159 243
rect 159 242 160 243
rect 160 242 161 243
rect 161 242 162 243
rect 162 242 163 243
rect 163 242 164 243
rect 164 242 165 243
rect 165 242 166 243
rect 166 242 167 243
rect 167 242 168 243
rect 168 242 169 243
rect 169 242 170 243
rect 170 242 171 243
rect 171 242 172 243
rect 172 242 173 243
rect 173 242 174 243
rect 174 242 175 243
rect 175 242 176 243
rect 176 242 177 243
rect 177 242 178 243
rect 178 242 179 243
rect 179 242 180 243
rect 180 242 181 243
rect 181 242 182 243
rect 182 242 183 243
rect 183 242 184 243
rect 184 242 185 243
rect 185 242 186 243
rect 186 242 187 243
rect 187 242 188 243
rect 214 242 215 243
rect 215 242 216 243
rect 216 242 217 243
rect 217 242 218 243
rect 218 242 219 243
rect 219 242 220 243
rect 220 242 221 243
rect 221 242 222 243
rect 222 242 223 243
rect 223 242 224 243
rect 224 242 225 243
rect 225 242 226 243
rect 226 242 227 243
rect 227 242 228 243
rect 228 242 229 243
rect 229 242 230 243
rect 230 242 231 243
rect 231 242 232 243
rect 232 242 233 243
rect 233 242 234 243
rect 234 242 235 243
rect 235 242 236 243
rect 236 242 237 243
rect 237 242 238 243
rect 238 242 239 243
rect 239 242 240 243
rect 240 242 241 243
rect 241 242 242 243
rect 242 242 243 243
rect 243 242 244 243
rect 246 242 247 243
rect 247 242 248 243
rect 248 242 249 243
rect 249 242 250 243
rect 250 242 251 243
rect 251 242 252 243
rect 252 242 253 243
rect 253 242 254 243
rect 254 242 255 243
rect 255 242 256 243
rect 257 242 258 243
rect 258 242 259 243
rect 259 242 260 243
rect 260 242 261 243
rect 261 242 262 243
rect 262 242 263 243
rect 263 242 264 243
rect 264 242 265 243
rect 265 242 266 243
rect 266 242 267 243
rect 267 242 268 243
rect 268 242 269 243
rect 269 242 270 243
rect 270 242 271 243
rect 271 242 272 243
rect 272 242 273 243
rect 273 242 274 243
rect 274 242 275 243
rect 275 242 276 243
rect 276 242 277 243
rect 277 242 278 243
rect 278 242 279 243
rect 279 242 280 243
rect 280 242 281 243
rect 281 242 282 243
rect 282 242 283 243
rect 283 242 284 243
rect 284 242 285 243
rect 285 242 286 243
rect 286 242 287 243
rect 287 242 288 243
rect 288 242 289 243
rect 315 242 316 243
rect 316 242 317 243
rect 317 242 318 243
rect 318 242 319 243
rect 372 242 373 243
rect 373 242 374 243
rect 374 242 375 243
rect 375 242 376 243
rect 376 242 377 243
rect 377 242 378 243
rect 378 242 379 243
rect 379 242 380 243
rect 380 242 381 243
rect 381 242 382 243
rect 382 242 383 243
rect 383 242 384 243
rect 384 242 385 243
rect 385 242 386 243
rect 386 242 387 243
rect 387 242 388 243
rect 388 242 389 243
rect 389 242 390 243
rect 390 242 391 243
rect 391 242 392 243
rect 392 242 393 243
rect 393 242 394 243
rect 394 242 395 243
rect 395 242 396 243
rect 396 242 397 243
rect 397 242 398 243
rect 398 242 399 243
rect 399 242 400 243
rect 74 241 75 242
rect 75 241 76 242
rect 76 241 77 242
rect 77 241 78 242
rect 78 241 79 242
rect 79 241 80 242
rect 80 241 81 242
rect 81 241 82 242
rect 82 241 83 242
rect 83 241 84 242
rect 84 241 85 242
rect 85 241 86 242
rect 86 241 87 242
rect 87 241 88 242
rect 97 241 98 242
rect 98 241 99 242
rect 99 241 100 242
rect 100 241 101 242
rect 101 241 102 242
rect 102 241 103 242
rect 103 241 104 242
rect 113 241 114 242
rect 114 241 115 242
rect 115 241 116 242
rect 116 241 117 242
rect 117 241 118 242
rect 118 241 119 242
rect 119 241 120 242
rect 120 241 121 242
rect 121 241 122 242
rect 122 241 123 242
rect 123 241 124 242
rect 124 241 125 242
rect 125 241 126 242
rect 126 241 127 242
rect 127 241 128 242
rect 128 241 129 242
rect 129 241 130 242
rect 130 241 131 242
rect 131 241 132 242
rect 132 241 133 242
rect 133 241 134 242
rect 134 241 135 242
rect 135 241 136 242
rect 136 241 137 242
rect 137 241 138 242
rect 138 241 139 242
rect 139 241 140 242
rect 140 241 141 242
rect 141 241 142 242
rect 142 241 143 242
rect 143 241 144 242
rect 144 241 145 242
rect 145 241 146 242
rect 146 241 147 242
rect 147 241 148 242
rect 148 241 149 242
rect 149 241 150 242
rect 150 241 151 242
rect 151 241 152 242
rect 152 241 153 242
rect 153 241 154 242
rect 154 241 155 242
rect 155 241 156 242
rect 156 241 157 242
rect 157 241 158 242
rect 158 241 159 242
rect 159 241 160 242
rect 160 241 161 242
rect 161 241 162 242
rect 162 241 163 242
rect 163 241 164 242
rect 164 241 165 242
rect 165 241 166 242
rect 166 241 167 242
rect 167 241 168 242
rect 168 241 169 242
rect 169 241 170 242
rect 170 241 171 242
rect 171 241 172 242
rect 172 241 173 242
rect 173 241 174 242
rect 174 241 175 242
rect 175 241 176 242
rect 176 241 177 242
rect 177 241 178 242
rect 178 241 179 242
rect 179 241 180 242
rect 180 241 181 242
rect 181 241 182 242
rect 182 241 183 242
rect 183 241 184 242
rect 184 241 185 242
rect 185 241 186 242
rect 186 241 187 242
rect 187 241 188 242
rect 188 241 189 242
rect 213 241 214 242
rect 214 241 215 242
rect 215 241 216 242
rect 216 241 217 242
rect 217 241 218 242
rect 218 241 219 242
rect 219 241 220 242
rect 220 241 221 242
rect 221 241 222 242
rect 222 241 223 242
rect 223 241 224 242
rect 224 241 225 242
rect 225 241 226 242
rect 226 241 227 242
rect 227 241 228 242
rect 228 241 229 242
rect 229 241 230 242
rect 230 241 231 242
rect 231 241 232 242
rect 232 241 233 242
rect 233 241 234 242
rect 234 241 235 242
rect 235 241 236 242
rect 236 241 237 242
rect 237 241 238 242
rect 238 241 239 242
rect 239 241 240 242
rect 240 241 241 242
rect 241 241 242 242
rect 242 241 243 242
rect 243 241 244 242
rect 244 241 245 242
rect 247 241 248 242
rect 248 241 249 242
rect 249 241 250 242
rect 250 241 251 242
rect 251 241 252 242
rect 252 241 253 242
rect 253 241 254 242
rect 254 241 255 242
rect 255 241 256 242
rect 256 241 257 242
rect 258 241 259 242
rect 259 241 260 242
rect 260 241 261 242
rect 261 241 262 242
rect 262 241 263 242
rect 263 241 264 242
rect 264 241 265 242
rect 265 241 266 242
rect 266 241 267 242
rect 267 241 268 242
rect 268 241 269 242
rect 269 241 270 242
rect 270 241 271 242
rect 271 241 272 242
rect 272 241 273 242
rect 273 241 274 242
rect 274 241 275 242
rect 275 241 276 242
rect 276 241 277 242
rect 277 241 278 242
rect 278 241 279 242
rect 279 241 280 242
rect 280 241 281 242
rect 281 241 282 242
rect 282 241 283 242
rect 283 241 284 242
rect 284 241 285 242
rect 285 241 286 242
rect 286 241 287 242
rect 287 241 288 242
rect 317 241 318 242
rect 318 241 319 242
rect 371 241 372 242
rect 372 241 373 242
rect 373 241 374 242
rect 374 241 375 242
rect 375 241 376 242
rect 376 241 377 242
rect 377 241 378 242
rect 378 241 379 242
rect 379 241 380 242
rect 383 241 384 242
rect 384 241 385 242
rect 385 241 386 242
rect 386 241 387 242
rect 387 241 388 242
rect 388 241 389 242
rect 389 241 390 242
rect 390 241 391 242
rect 391 241 392 242
rect 392 241 393 242
rect 393 241 394 242
rect 394 241 395 242
rect 395 241 396 242
rect 396 241 397 242
rect 397 241 398 242
rect 398 241 399 242
rect 399 241 400 242
rect 400 241 401 242
rect 401 241 402 242
rect 402 241 403 242
rect 403 241 404 242
rect 75 240 76 241
rect 76 240 77 241
rect 77 240 78 241
rect 78 240 79 241
rect 79 240 80 241
rect 80 240 81 241
rect 81 240 82 241
rect 82 240 83 241
rect 83 240 84 241
rect 84 240 85 241
rect 85 240 86 241
rect 86 240 87 241
rect 87 240 88 241
rect 88 240 89 241
rect 89 240 90 241
rect 98 240 99 241
rect 99 240 100 241
rect 100 240 101 241
rect 101 240 102 241
rect 102 240 103 241
rect 103 240 104 241
rect 104 240 105 241
rect 105 240 106 241
rect 106 240 107 241
rect 107 240 108 241
rect 108 240 109 241
rect 109 240 110 241
rect 110 240 111 241
rect 111 240 112 241
rect 112 240 113 241
rect 113 240 114 241
rect 114 240 115 241
rect 115 240 116 241
rect 116 240 117 241
rect 117 240 118 241
rect 118 240 119 241
rect 119 240 120 241
rect 120 240 121 241
rect 121 240 122 241
rect 122 240 123 241
rect 123 240 124 241
rect 124 240 125 241
rect 125 240 126 241
rect 126 240 127 241
rect 127 240 128 241
rect 128 240 129 241
rect 129 240 130 241
rect 130 240 131 241
rect 131 240 132 241
rect 132 240 133 241
rect 133 240 134 241
rect 134 240 135 241
rect 135 240 136 241
rect 136 240 137 241
rect 137 240 138 241
rect 138 240 139 241
rect 139 240 140 241
rect 140 240 141 241
rect 141 240 142 241
rect 142 240 143 241
rect 143 240 144 241
rect 144 240 145 241
rect 145 240 146 241
rect 146 240 147 241
rect 147 240 148 241
rect 148 240 149 241
rect 149 240 150 241
rect 150 240 151 241
rect 151 240 152 241
rect 152 240 153 241
rect 153 240 154 241
rect 154 240 155 241
rect 155 240 156 241
rect 156 240 157 241
rect 157 240 158 241
rect 158 240 159 241
rect 159 240 160 241
rect 160 240 161 241
rect 161 240 162 241
rect 162 240 163 241
rect 163 240 164 241
rect 164 240 165 241
rect 165 240 166 241
rect 166 240 167 241
rect 167 240 168 241
rect 168 240 169 241
rect 169 240 170 241
rect 170 240 171 241
rect 171 240 172 241
rect 172 240 173 241
rect 173 240 174 241
rect 174 240 175 241
rect 175 240 176 241
rect 176 240 177 241
rect 177 240 178 241
rect 178 240 179 241
rect 179 240 180 241
rect 180 240 181 241
rect 181 240 182 241
rect 182 240 183 241
rect 183 240 184 241
rect 184 240 185 241
rect 185 240 186 241
rect 186 240 187 241
rect 187 240 188 241
rect 188 240 189 241
rect 213 240 214 241
rect 214 240 215 241
rect 215 240 216 241
rect 216 240 217 241
rect 217 240 218 241
rect 218 240 219 241
rect 219 240 220 241
rect 220 240 221 241
rect 221 240 222 241
rect 222 240 223 241
rect 223 240 224 241
rect 224 240 225 241
rect 225 240 226 241
rect 226 240 227 241
rect 227 240 228 241
rect 228 240 229 241
rect 229 240 230 241
rect 230 240 231 241
rect 231 240 232 241
rect 232 240 233 241
rect 233 240 234 241
rect 234 240 235 241
rect 235 240 236 241
rect 236 240 237 241
rect 237 240 238 241
rect 238 240 239 241
rect 239 240 240 241
rect 240 240 241 241
rect 241 240 242 241
rect 242 240 243 241
rect 243 240 244 241
rect 244 240 245 241
rect 245 240 246 241
rect 246 240 247 241
rect 248 240 249 241
rect 249 240 250 241
rect 250 240 251 241
rect 251 240 252 241
rect 252 240 253 241
rect 253 240 254 241
rect 254 240 255 241
rect 255 240 256 241
rect 256 240 257 241
rect 257 240 258 241
rect 258 240 259 241
rect 259 240 260 241
rect 260 240 261 241
rect 261 240 262 241
rect 262 240 263 241
rect 263 240 264 241
rect 264 240 265 241
rect 265 240 266 241
rect 266 240 267 241
rect 267 240 268 241
rect 268 240 269 241
rect 269 240 270 241
rect 270 240 271 241
rect 271 240 272 241
rect 272 240 273 241
rect 273 240 274 241
rect 274 240 275 241
rect 275 240 276 241
rect 276 240 277 241
rect 277 240 278 241
rect 278 240 279 241
rect 279 240 280 241
rect 280 240 281 241
rect 281 240 282 241
rect 282 240 283 241
rect 283 240 284 241
rect 284 240 285 241
rect 285 240 286 241
rect 335 240 336 241
rect 370 240 371 241
rect 371 240 372 241
rect 372 240 373 241
rect 373 240 374 241
rect 374 240 375 241
rect 375 240 376 241
rect 376 240 377 241
rect 377 240 378 241
rect 378 240 379 241
rect 385 240 386 241
rect 386 240 387 241
rect 387 240 388 241
rect 388 240 389 241
rect 389 240 390 241
rect 390 240 391 241
rect 391 240 392 241
rect 392 240 393 241
rect 393 240 394 241
rect 394 240 395 241
rect 395 240 396 241
rect 396 240 397 241
rect 397 240 398 241
rect 398 240 399 241
rect 399 240 400 241
rect 400 240 401 241
rect 401 240 402 241
rect 402 240 403 241
rect 403 240 404 241
rect 404 240 405 241
rect 405 240 406 241
rect 406 240 407 241
rect 407 240 408 241
rect 408 240 409 241
rect 77 239 78 240
rect 78 239 79 240
rect 79 239 80 240
rect 80 239 81 240
rect 81 239 82 240
rect 82 239 83 240
rect 83 239 84 240
rect 84 239 85 240
rect 85 239 86 240
rect 86 239 87 240
rect 87 239 88 240
rect 88 239 89 240
rect 89 239 90 240
rect 90 239 91 240
rect 100 239 101 240
rect 101 239 102 240
rect 102 239 103 240
rect 103 239 104 240
rect 104 239 105 240
rect 105 239 106 240
rect 106 239 107 240
rect 107 239 108 240
rect 108 239 109 240
rect 109 239 110 240
rect 110 239 111 240
rect 111 239 112 240
rect 112 239 113 240
rect 113 239 114 240
rect 114 239 115 240
rect 115 239 116 240
rect 116 239 117 240
rect 117 239 118 240
rect 118 239 119 240
rect 119 239 120 240
rect 120 239 121 240
rect 121 239 122 240
rect 122 239 123 240
rect 123 239 124 240
rect 124 239 125 240
rect 125 239 126 240
rect 126 239 127 240
rect 127 239 128 240
rect 128 239 129 240
rect 129 239 130 240
rect 130 239 131 240
rect 131 239 132 240
rect 132 239 133 240
rect 133 239 134 240
rect 134 239 135 240
rect 135 239 136 240
rect 136 239 137 240
rect 137 239 138 240
rect 138 239 139 240
rect 139 239 140 240
rect 140 239 141 240
rect 141 239 142 240
rect 142 239 143 240
rect 143 239 144 240
rect 144 239 145 240
rect 145 239 146 240
rect 146 239 147 240
rect 147 239 148 240
rect 148 239 149 240
rect 149 239 150 240
rect 150 239 151 240
rect 151 239 152 240
rect 152 239 153 240
rect 153 239 154 240
rect 154 239 155 240
rect 155 239 156 240
rect 156 239 157 240
rect 157 239 158 240
rect 158 239 159 240
rect 159 239 160 240
rect 160 239 161 240
rect 161 239 162 240
rect 162 239 163 240
rect 163 239 164 240
rect 164 239 165 240
rect 165 239 166 240
rect 166 239 167 240
rect 167 239 168 240
rect 168 239 169 240
rect 169 239 170 240
rect 170 239 171 240
rect 171 239 172 240
rect 172 239 173 240
rect 173 239 174 240
rect 174 239 175 240
rect 175 239 176 240
rect 176 239 177 240
rect 177 239 178 240
rect 178 239 179 240
rect 179 239 180 240
rect 180 239 181 240
rect 181 239 182 240
rect 183 239 184 240
rect 184 239 185 240
rect 185 239 186 240
rect 186 239 187 240
rect 187 239 188 240
rect 188 239 189 240
rect 212 239 213 240
rect 213 239 214 240
rect 214 239 215 240
rect 215 239 216 240
rect 216 239 217 240
rect 217 239 218 240
rect 218 239 219 240
rect 219 239 220 240
rect 220 239 221 240
rect 221 239 222 240
rect 222 239 223 240
rect 223 239 224 240
rect 224 239 225 240
rect 225 239 226 240
rect 226 239 227 240
rect 227 239 228 240
rect 228 239 229 240
rect 229 239 230 240
rect 230 239 231 240
rect 231 239 232 240
rect 232 239 233 240
rect 233 239 234 240
rect 234 239 235 240
rect 235 239 236 240
rect 236 239 237 240
rect 237 239 238 240
rect 238 239 239 240
rect 239 239 240 240
rect 240 239 241 240
rect 241 239 242 240
rect 242 239 243 240
rect 243 239 244 240
rect 244 239 245 240
rect 245 239 246 240
rect 246 239 247 240
rect 247 239 248 240
rect 250 239 251 240
rect 251 239 252 240
rect 252 239 253 240
rect 253 239 254 240
rect 254 239 255 240
rect 255 239 256 240
rect 256 239 257 240
rect 257 239 258 240
rect 258 239 259 240
rect 259 239 260 240
rect 260 239 261 240
rect 261 239 262 240
rect 262 239 263 240
rect 263 239 264 240
rect 264 239 265 240
rect 265 239 266 240
rect 266 239 267 240
rect 267 239 268 240
rect 268 239 269 240
rect 269 239 270 240
rect 270 239 271 240
rect 271 239 272 240
rect 272 239 273 240
rect 273 239 274 240
rect 274 239 275 240
rect 275 239 276 240
rect 276 239 277 240
rect 277 239 278 240
rect 278 239 279 240
rect 279 239 280 240
rect 280 239 281 240
rect 281 239 282 240
rect 282 239 283 240
rect 283 239 284 240
rect 284 239 285 240
rect 335 239 336 240
rect 369 239 370 240
rect 370 239 371 240
rect 371 239 372 240
rect 372 239 373 240
rect 373 239 374 240
rect 374 239 375 240
rect 375 239 376 240
rect 376 239 377 240
rect 377 239 378 240
rect 388 239 389 240
rect 389 239 390 240
rect 390 239 391 240
rect 391 239 392 240
rect 392 239 393 240
rect 393 239 394 240
rect 394 239 395 240
rect 395 239 396 240
rect 396 239 397 240
rect 397 239 398 240
rect 398 239 399 240
rect 399 239 400 240
rect 400 239 401 240
rect 401 239 402 240
rect 402 239 403 240
rect 403 239 404 240
rect 404 239 405 240
rect 405 239 406 240
rect 406 239 407 240
rect 407 239 408 240
rect 408 239 409 240
rect 409 239 410 240
rect 410 239 411 240
rect 411 239 412 240
rect 78 238 79 239
rect 79 238 80 239
rect 80 238 81 239
rect 81 238 82 239
rect 82 238 83 239
rect 83 238 84 239
rect 84 238 85 239
rect 85 238 86 239
rect 86 238 87 239
rect 87 238 88 239
rect 88 238 89 239
rect 89 238 90 239
rect 90 238 91 239
rect 91 238 92 239
rect 92 238 93 239
rect 101 238 102 239
rect 102 238 103 239
rect 103 238 104 239
rect 104 238 105 239
rect 105 238 106 239
rect 106 238 107 239
rect 107 238 108 239
rect 108 238 109 239
rect 109 238 110 239
rect 110 238 111 239
rect 111 238 112 239
rect 112 238 113 239
rect 113 238 114 239
rect 114 238 115 239
rect 115 238 116 239
rect 116 238 117 239
rect 117 238 118 239
rect 118 238 119 239
rect 119 238 120 239
rect 120 238 121 239
rect 121 238 122 239
rect 122 238 123 239
rect 123 238 124 239
rect 124 238 125 239
rect 125 238 126 239
rect 126 238 127 239
rect 127 238 128 239
rect 128 238 129 239
rect 129 238 130 239
rect 130 238 131 239
rect 131 238 132 239
rect 132 238 133 239
rect 133 238 134 239
rect 134 238 135 239
rect 135 238 136 239
rect 136 238 137 239
rect 137 238 138 239
rect 138 238 139 239
rect 139 238 140 239
rect 140 238 141 239
rect 141 238 142 239
rect 142 238 143 239
rect 143 238 144 239
rect 144 238 145 239
rect 145 238 146 239
rect 146 238 147 239
rect 147 238 148 239
rect 148 238 149 239
rect 149 238 150 239
rect 150 238 151 239
rect 151 238 152 239
rect 152 238 153 239
rect 153 238 154 239
rect 154 238 155 239
rect 155 238 156 239
rect 156 238 157 239
rect 157 238 158 239
rect 158 238 159 239
rect 159 238 160 239
rect 160 238 161 239
rect 161 238 162 239
rect 162 238 163 239
rect 163 238 164 239
rect 164 238 165 239
rect 165 238 166 239
rect 166 238 167 239
rect 167 238 168 239
rect 168 238 169 239
rect 169 238 170 239
rect 170 238 171 239
rect 171 238 172 239
rect 172 238 173 239
rect 173 238 174 239
rect 174 238 175 239
rect 175 238 176 239
rect 176 238 177 239
rect 177 238 178 239
rect 178 238 179 239
rect 179 238 180 239
rect 184 238 185 239
rect 185 238 186 239
rect 186 238 187 239
rect 187 238 188 239
rect 188 238 189 239
rect 189 238 190 239
rect 211 238 212 239
rect 212 238 213 239
rect 213 238 214 239
rect 214 238 215 239
rect 215 238 216 239
rect 216 238 217 239
rect 217 238 218 239
rect 218 238 219 239
rect 219 238 220 239
rect 220 238 221 239
rect 221 238 222 239
rect 222 238 223 239
rect 223 238 224 239
rect 224 238 225 239
rect 225 238 226 239
rect 226 238 227 239
rect 227 238 228 239
rect 228 238 229 239
rect 229 238 230 239
rect 230 238 231 239
rect 231 238 232 239
rect 232 238 233 239
rect 233 238 234 239
rect 234 238 235 239
rect 235 238 236 239
rect 236 238 237 239
rect 237 238 238 239
rect 238 238 239 239
rect 239 238 240 239
rect 240 238 241 239
rect 241 238 242 239
rect 242 238 243 239
rect 243 238 244 239
rect 244 238 245 239
rect 245 238 246 239
rect 246 238 247 239
rect 247 238 248 239
rect 248 238 249 239
rect 249 238 250 239
rect 251 238 252 239
rect 252 238 253 239
rect 253 238 254 239
rect 254 238 255 239
rect 255 238 256 239
rect 256 238 257 239
rect 257 238 258 239
rect 258 238 259 239
rect 259 238 260 239
rect 260 238 261 239
rect 261 238 262 239
rect 262 238 263 239
rect 263 238 264 239
rect 264 238 265 239
rect 265 238 266 239
rect 266 238 267 239
rect 267 238 268 239
rect 268 238 269 239
rect 269 238 270 239
rect 270 238 271 239
rect 271 238 272 239
rect 272 238 273 239
rect 273 238 274 239
rect 274 238 275 239
rect 275 238 276 239
rect 276 238 277 239
rect 277 238 278 239
rect 278 238 279 239
rect 279 238 280 239
rect 280 238 281 239
rect 281 238 282 239
rect 282 238 283 239
rect 283 238 284 239
rect 335 238 336 239
rect 336 238 337 239
rect 368 238 369 239
rect 369 238 370 239
rect 370 238 371 239
rect 371 238 372 239
rect 372 238 373 239
rect 373 238 374 239
rect 374 238 375 239
rect 375 238 376 239
rect 376 238 377 239
rect 391 238 392 239
rect 392 238 393 239
rect 393 238 394 239
rect 394 238 395 239
rect 395 238 396 239
rect 396 238 397 239
rect 397 238 398 239
rect 398 238 399 239
rect 399 238 400 239
rect 400 238 401 239
rect 401 238 402 239
rect 402 238 403 239
rect 403 238 404 239
rect 404 238 405 239
rect 405 238 406 239
rect 406 238 407 239
rect 407 238 408 239
rect 408 238 409 239
rect 409 238 410 239
rect 410 238 411 239
rect 79 237 80 238
rect 80 237 81 238
rect 81 237 82 238
rect 82 237 83 238
rect 83 237 84 238
rect 84 237 85 238
rect 85 237 86 238
rect 86 237 87 238
rect 87 237 88 238
rect 88 237 89 238
rect 89 237 90 238
rect 90 237 91 238
rect 91 237 92 238
rect 92 237 93 238
rect 93 237 94 238
rect 102 237 103 238
rect 103 237 104 238
rect 104 237 105 238
rect 105 237 106 238
rect 106 237 107 238
rect 107 237 108 238
rect 108 237 109 238
rect 109 237 110 238
rect 110 237 111 238
rect 111 237 112 238
rect 112 237 113 238
rect 113 237 114 238
rect 114 237 115 238
rect 115 237 116 238
rect 116 237 117 238
rect 117 237 118 238
rect 118 237 119 238
rect 119 237 120 238
rect 120 237 121 238
rect 121 237 122 238
rect 122 237 123 238
rect 123 237 124 238
rect 124 237 125 238
rect 125 237 126 238
rect 126 237 127 238
rect 127 237 128 238
rect 128 237 129 238
rect 129 237 130 238
rect 130 237 131 238
rect 131 237 132 238
rect 132 237 133 238
rect 133 237 134 238
rect 134 237 135 238
rect 135 237 136 238
rect 136 237 137 238
rect 137 237 138 238
rect 138 237 139 238
rect 139 237 140 238
rect 140 237 141 238
rect 141 237 142 238
rect 142 237 143 238
rect 143 237 144 238
rect 144 237 145 238
rect 145 237 146 238
rect 146 237 147 238
rect 147 237 148 238
rect 148 237 149 238
rect 149 237 150 238
rect 150 237 151 238
rect 151 237 152 238
rect 152 237 153 238
rect 153 237 154 238
rect 154 237 155 238
rect 155 237 156 238
rect 156 237 157 238
rect 157 237 158 238
rect 158 237 159 238
rect 159 237 160 238
rect 160 237 161 238
rect 161 237 162 238
rect 162 237 163 238
rect 163 237 164 238
rect 164 237 165 238
rect 165 237 166 238
rect 166 237 167 238
rect 167 237 168 238
rect 168 237 169 238
rect 169 237 170 238
rect 170 237 171 238
rect 171 237 172 238
rect 172 237 173 238
rect 173 237 174 238
rect 174 237 175 238
rect 175 237 176 238
rect 176 237 177 238
rect 177 237 178 238
rect 178 237 179 238
rect 184 237 185 238
rect 185 237 186 238
rect 186 237 187 238
rect 187 237 188 238
rect 188 237 189 238
rect 189 237 190 238
rect 190 237 191 238
rect 210 237 211 238
rect 211 237 212 238
rect 212 237 213 238
rect 213 237 214 238
rect 214 237 215 238
rect 215 237 216 238
rect 216 237 217 238
rect 217 237 218 238
rect 218 237 219 238
rect 219 237 220 238
rect 220 237 221 238
rect 221 237 222 238
rect 222 237 223 238
rect 223 237 224 238
rect 224 237 225 238
rect 225 237 226 238
rect 226 237 227 238
rect 227 237 228 238
rect 228 237 229 238
rect 229 237 230 238
rect 230 237 231 238
rect 231 237 232 238
rect 232 237 233 238
rect 233 237 234 238
rect 234 237 235 238
rect 235 237 236 238
rect 236 237 237 238
rect 237 237 238 238
rect 238 237 239 238
rect 239 237 240 238
rect 240 237 241 238
rect 241 237 242 238
rect 242 237 243 238
rect 243 237 244 238
rect 244 237 245 238
rect 245 237 246 238
rect 246 237 247 238
rect 247 237 248 238
rect 248 237 249 238
rect 249 237 250 238
rect 250 237 251 238
rect 251 237 252 238
rect 252 237 253 238
rect 253 237 254 238
rect 254 237 255 238
rect 255 237 256 238
rect 256 237 257 238
rect 257 237 258 238
rect 258 237 259 238
rect 259 237 260 238
rect 260 237 261 238
rect 261 237 262 238
rect 262 237 263 238
rect 263 237 264 238
rect 264 237 265 238
rect 265 237 266 238
rect 266 237 267 238
rect 267 237 268 238
rect 268 237 269 238
rect 269 237 270 238
rect 270 237 271 238
rect 271 237 272 238
rect 272 237 273 238
rect 273 237 274 238
rect 274 237 275 238
rect 275 237 276 238
rect 276 237 277 238
rect 277 237 278 238
rect 278 237 279 238
rect 279 237 280 238
rect 280 237 281 238
rect 281 237 282 238
rect 335 237 336 238
rect 336 237 337 238
rect 367 237 368 238
rect 368 237 369 238
rect 369 237 370 238
rect 370 237 371 238
rect 371 237 372 238
rect 372 237 373 238
rect 373 237 374 238
rect 374 237 375 238
rect 375 237 376 238
rect 376 237 377 238
rect 394 237 395 238
rect 395 237 396 238
rect 396 237 397 238
rect 397 237 398 238
rect 398 237 399 238
rect 399 237 400 238
rect 400 237 401 238
rect 401 237 402 238
rect 402 237 403 238
rect 403 237 404 238
rect 404 237 405 238
rect 405 237 406 238
rect 406 237 407 238
rect 407 237 408 238
rect 408 237 409 238
rect 409 237 410 238
rect 410 237 411 238
rect 80 236 81 237
rect 81 236 82 237
rect 82 236 83 237
rect 83 236 84 237
rect 84 236 85 237
rect 85 236 86 237
rect 86 236 87 237
rect 87 236 88 237
rect 88 236 89 237
rect 89 236 90 237
rect 90 236 91 237
rect 91 236 92 237
rect 92 236 93 237
rect 93 236 94 237
rect 94 236 95 237
rect 95 236 96 237
rect 104 236 105 237
rect 105 236 106 237
rect 106 236 107 237
rect 107 236 108 237
rect 108 236 109 237
rect 109 236 110 237
rect 110 236 111 237
rect 111 236 112 237
rect 112 236 113 237
rect 113 236 114 237
rect 114 236 115 237
rect 115 236 116 237
rect 116 236 117 237
rect 117 236 118 237
rect 118 236 119 237
rect 119 236 120 237
rect 120 236 121 237
rect 121 236 122 237
rect 122 236 123 237
rect 123 236 124 237
rect 124 236 125 237
rect 125 236 126 237
rect 126 236 127 237
rect 127 236 128 237
rect 128 236 129 237
rect 129 236 130 237
rect 130 236 131 237
rect 131 236 132 237
rect 132 236 133 237
rect 133 236 134 237
rect 134 236 135 237
rect 135 236 136 237
rect 136 236 137 237
rect 137 236 138 237
rect 138 236 139 237
rect 139 236 140 237
rect 140 236 141 237
rect 141 236 142 237
rect 142 236 143 237
rect 143 236 144 237
rect 144 236 145 237
rect 145 236 146 237
rect 146 236 147 237
rect 147 236 148 237
rect 148 236 149 237
rect 149 236 150 237
rect 150 236 151 237
rect 151 236 152 237
rect 152 236 153 237
rect 153 236 154 237
rect 154 236 155 237
rect 155 236 156 237
rect 156 236 157 237
rect 157 236 158 237
rect 158 236 159 237
rect 159 236 160 237
rect 160 236 161 237
rect 161 236 162 237
rect 162 236 163 237
rect 163 236 164 237
rect 164 236 165 237
rect 165 236 166 237
rect 166 236 167 237
rect 167 236 168 237
rect 168 236 169 237
rect 169 236 170 237
rect 170 236 171 237
rect 171 236 172 237
rect 172 236 173 237
rect 173 236 174 237
rect 174 236 175 237
rect 175 236 176 237
rect 176 236 177 237
rect 184 236 185 237
rect 185 236 186 237
rect 186 236 187 237
rect 187 236 188 237
rect 188 236 189 237
rect 189 236 190 237
rect 190 236 191 237
rect 191 236 192 237
rect 209 236 210 237
rect 210 236 211 237
rect 211 236 212 237
rect 212 236 213 237
rect 213 236 214 237
rect 214 236 215 237
rect 215 236 216 237
rect 221 236 222 237
rect 222 236 223 237
rect 223 236 224 237
rect 224 236 225 237
rect 225 236 226 237
rect 226 236 227 237
rect 227 236 228 237
rect 228 236 229 237
rect 229 236 230 237
rect 230 236 231 237
rect 231 236 232 237
rect 232 236 233 237
rect 233 236 234 237
rect 234 236 235 237
rect 235 236 236 237
rect 236 236 237 237
rect 237 236 238 237
rect 238 236 239 237
rect 239 236 240 237
rect 240 236 241 237
rect 241 236 242 237
rect 242 236 243 237
rect 243 236 244 237
rect 244 236 245 237
rect 245 236 246 237
rect 246 236 247 237
rect 247 236 248 237
rect 248 236 249 237
rect 249 236 250 237
rect 250 236 251 237
rect 251 236 252 237
rect 252 236 253 237
rect 253 236 254 237
rect 254 236 255 237
rect 255 236 256 237
rect 256 236 257 237
rect 257 236 258 237
rect 258 236 259 237
rect 259 236 260 237
rect 260 236 261 237
rect 261 236 262 237
rect 262 236 263 237
rect 263 236 264 237
rect 264 236 265 237
rect 265 236 266 237
rect 266 236 267 237
rect 267 236 268 237
rect 268 236 269 237
rect 269 236 270 237
rect 270 236 271 237
rect 271 236 272 237
rect 272 236 273 237
rect 273 236 274 237
rect 274 236 275 237
rect 275 236 276 237
rect 276 236 277 237
rect 277 236 278 237
rect 278 236 279 237
rect 279 236 280 237
rect 335 236 336 237
rect 336 236 337 237
rect 366 236 367 237
rect 367 236 368 237
rect 368 236 369 237
rect 369 236 370 237
rect 370 236 371 237
rect 371 236 372 237
rect 372 236 373 237
rect 373 236 374 237
rect 374 236 375 237
rect 375 236 376 237
rect 398 236 399 237
rect 399 236 400 237
rect 400 236 401 237
rect 401 236 402 237
rect 402 236 403 237
rect 403 236 404 237
rect 404 236 405 237
rect 405 236 406 237
rect 406 236 407 237
rect 407 236 408 237
rect 408 236 409 237
rect 409 236 410 237
rect 81 235 82 236
rect 82 235 83 236
rect 83 235 84 236
rect 84 235 85 236
rect 85 235 86 236
rect 86 235 87 236
rect 87 235 88 236
rect 88 235 89 236
rect 89 235 90 236
rect 90 235 91 236
rect 91 235 92 236
rect 92 235 93 236
rect 93 235 94 236
rect 94 235 95 236
rect 95 235 96 236
rect 96 235 97 236
rect 97 235 98 236
rect 106 235 107 236
rect 107 235 108 236
rect 108 235 109 236
rect 109 235 110 236
rect 110 235 111 236
rect 111 235 112 236
rect 112 235 113 236
rect 113 235 114 236
rect 114 235 115 236
rect 115 235 116 236
rect 116 235 117 236
rect 117 235 118 236
rect 118 235 119 236
rect 119 235 120 236
rect 120 235 121 236
rect 121 235 122 236
rect 122 235 123 236
rect 123 235 124 236
rect 124 235 125 236
rect 125 235 126 236
rect 126 235 127 236
rect 127 235 128 236
rect 128 235 129 236
rect 129 235 130 236
rect 130 235 131 236
rect 131 235 132 236
rect 132 235 133 236
rect 133 235 134 236
rect 134 235 135 236
rect 135 235 136 236
rect 136 235 137 236
rect 137 235 138 236
rect 138 235 139 236
rect 139 235 140 236
rect 140 235 141 236
rect 141 235 142 236
rect 142 235 143 236
rect 143 235 144 236
rect 144 235 145 236
rect 145 235 146 236
rect 146 235 147 236
rect 147 235 148 236
rect 148 235 149 236
rect 149 235 150 236
rect 150 235 151 236
rect 151 235 152 236
rect 152 235 153 236
rect 153 235 154 236
rect 154 235 155 236
rect 155 235 156 236
rect 156 235 157 236
rect 157 235 158 236
rect 158 235 159 236
rect 159 235 160 236
rect 160 235 161 236
rect 161 235 162 236
rect 162 235 163 236
rect 163 235 164 236
rect 164 235 165 236
rect 165 235 166 236
rect 166 235 167 236
rect 167 235 168 236
rect 168 235 169 236
rect 169 235 170 236
rect 170 235 171 236
rect 171 235 172 236
rect 172 235 173 236
rect 173 235 174 236
rect 174 235 175 236
rect 175 235 176 236
rect 185 235 186 236
rect 186 235 187 236
rect 187 235 188 236
rect 188 235 189 236
rect 189 235 190 236
rect 190 235 191 236
rect 191 235 192 236
rect 192 235 193 236
rect 208 235 209 236
rect 209 235 210 236
rect 210 235 211 236
rect 211 235 212 236
rect 212 235 213 236
rect 213 235 214 236
rect 214 235 215 236
rect 224 235 225 236
rect 225 235 226 236
rect 226 235 227 236
rect 227 235 228 236
rect 228 235 229 236
rect 229 235 230 236
rect 230 235 231 236
rect 231 235 232 236
rect 232 235 233 236
rect 233 235 234 236
rect 234 235 235 236
rect 235 235 236 236
rect 236 235 237 236
rect 237 235 238 236
rect 238 235 239 236
rect 239 235 240 236
rect 240 235 241 236
rect 241 235 242 236
rect 242 235 243 236
rect 243 235 244 236
rect 244 235 245 236
rect 245 235 246 236
rect 246 235 247 236
rect 247 235 248 236
rect 248 235 249 236
rect 249 235 250 236
rect 250 235 251 236
rect 251 235 252 236
rect 252 235 253 236
rect 253 235 254 236
rect 254 235 255 236
rect 255 235 256 236
rect 256 235 257 236
rect 257 235 258 236
rect 258 235 259 236
rect 259 235 260 236
rect 260 235 261 236
rect 261 235 262 236
rect 262 235 263 236
rect 263 235 264 236
rect 264 235 265 236
rect 265 235 266 236
rect 266 235 267 236
rect 267 235 268 236
rect 268 235 269 236
rect 269 235 270 236
rect 270 235 271 236
rect 271 235 272 236
rect 272 235 273 236
rect 273 235 274 236
rect 274 235 275 236
rect 275 235 276 236
rect 276 235 277 236
rect 277 235 278 236
rect 278 235 279 236
rect 334 235 335 236
rect 335 235 336 236
rect 336 235 337 236
rect 337 235 338 236
rect 365 235 366 236
rect 366 235 367 236
rect 367 235 368 236
rect 368 235 369 236
rect 369 235 370 236
rect 370 235 371 236
rect 371 235 372 236
rect 372 235 373 236
rect 373 235 374 236
rect 374 235 375 236
rect 402 235 403 236
rect 403 235 404 236
rect 404 235 405 236
rect 405 235 406 236
rect 406 235 407 236
rect 407 235 408 236
rect 408 235 409 236
rect 409 235 410 236
rect 83 234 84 235
rect 84 234 85 235
rect 85 234 86 235
rect 86 234 87 235
rect 87 234 88 235
rect 88 234 89 235
rect 89 234 90 235
rect 90 234 91 235
rect 91 234 92 235
rect 92 234 93 235
rect 93 234 94 235
rect 94 234 95 235
rect 95 234 96 235
rect 96 234 97 235
rect 97 234 98 235
rect 98 234 99 235
rect 107 234 108 235
rect 108 234 109 235
rect 109 234 110 235
rect 110 234 111 235
rect 111 234 112 235
rect 112 234 113 235
rect 113 234 114 235
rect 114 234 115 235
rect 115 234 116 235
rect 116 234 117 235
rect 117 234 118 235
rect 118 234 119 235
rect 119 234 120 235
rect 120 234 121 235
rect 121 234 122 235
rect 122 234 123 235
rect 123 234 124 235
rect 124 234 125 235
rect 125 234 126 235
rect 126 234 127 235
rect 127 234 128 235
rect 128 234 129 235
rect 129 234 130 235
rect 130 234 131 235
rect 131 234 132 235
rect 132 234 133 235
rect 133 234 134 235
rect 134 234 135 235
rect 135 234 136 235
rect 136 234 137 235
rect 137 234 138 235
rect 138 234 139 235
rect 139 234 140 235
rect 140 234 141 235
rect 141 234 142 235
rect 142 234 143 235
rect 143 234 144 235
rect 144 234 145 235
rect 145 234 146 235
rect 146 234 147 235
rect 147 234 148 235
rect 148 234 149 235
rect 149 234 150 235
rect 150 234 151 235
rect 151 234 152 235
rect 152 234 153 235
rect 153 234 154 235
rect 154 234 155 235
rect 155 234 156 235
rect 156 234 157 235
rect 157 234 158 235
rect 158 234 159 235
rect 159 234 160 235
rect 160 234 161 235
rect 161 234 162 235
rect 162 234 163 235
rect 163 234 164 235
rect 164 234 165 235
rect 165 234 166 235
rect 166 234 167 235
rect 167 234 168 235
rect 168 234 169 235
rect 169 234 170 235
rect 170 234 171 235
rect 171 234 172 235
rect 172 234 173 235
rect 173 234 174 235
rect 174 234 175 235
rect 185 234 186 235
rect 186 234 187 235
rect 187 234 188 235
rect 188 234 189 235
rect 189 234 190 235
rect 190 234 191 235
rect 191 234 192 235
rect 192 234 193 235
rect 193 234 194 235
rect 194 234 195 235
rect 206 234 207 235
rect 207 234 208 235
rect 208 234 209 235
rect 209 234 210 235
rect 210 234 211 235
rect 211 234 212 235
rect 212 234 213 235
rect 213 234 214 235
rect 214 234 215 235
rect 227 234 228 235
rect 228 234 229 235
rect 229 234 230 235
rect 230 234 231 235
rect 231 234 232 235
rect 232 234 233 235
rect 233 234 234 235
rect 234 234 235 235
rect 235 234 236 235
rect 236 234 237 235
rect 237 234 238 235
rect 238 234 239 235
rect 239 234 240 235
rect 240 234 241 235
rect 241 234 242 235
rect 242 234 243 235
rect 243 234 244 235
rect 244 234 245 235
rect 245 234 246 235
rect 246 234 247 235
rect 247 234 248 235
rect 248 234 249 235
rect 249 234 250 235
rect 250 234 251 235
rect 251 234 252 235
rect 252 234 253 235
rect 253 234 254 235
rect 254 234 255 235
rect 255 234 256 235
rect 256 234 257 235
rect 257 234 258 235
rect 258 234 259 235
rect 259 234 260 235
rect 260 234 261 235
rect 261 234 262 235
rect 262 234 263 235
rect 263 234 264 235
rect 264 234 265 235
rect 265 234 266 235
rect 266 234 267 235
rect 267 234 268 235
rect 268 234 269 235
rect 269 234 270 235
rect 270 234 271 235
rect 271 234 272 235
rect 272 234 273 235
rect 273 234 274 235
rect 274 234 275 235
rect 275 234 276 235
rect 276 234 277 235
rect 277 234 278 235
rect 278 234 279 235
rect 279 234 280 235
rect 280 234 281 235
rect 334 234 335 235
rect 335 234 336 235
rect 336 234 337 235
rect 337 234 338 235
rect 338 234 339 235
rect 364 234 365 235
rect 365 234 366 235
rect 366 234 367 235
rect 367 234 368 235
rect 368 234 369 235
rect 369 234 370 235
rect 370 234 371 235
rect 371 234 372 235
rect 372 234 373 235
rect 373 234 374 235
rect 402 234 403 235
rect 403 234 404 235
rect 404 234 405 235
rect 405 234 406 235
rect 406 234 407 235
rect 407 234 408 235
rect 408 234 409 235
rect 84 233 85 234
rect 85 233 86 234
rect 86 233 87 234
rect 87 233 88 234
rect 88 233 89 234
rect 89 233 90 234
rect 90 233 91 234
rect 91 233 92 234
rect 92 233 93 234
rect 93 233 94 234
rect 94 233 95 234
rect 95 233 96 234
rect 96 233 97 234
rect 97 233 98 234
rect 98 233 99 234
rect 99 233 100 234
rect 100 233 101 234
rect 101 233 102 234
rect 110 233 111 234
rect 111 233 112 234
rect 112 233 113 234
rect 113 233 114 234
rect 114 233 115 234
rect 115 233 116 234
rect 116 233 117 234
rect 117 233 118 234
rect 118 233 119 234
rect 119 233 120 234
rect 120 233 121 234
rect 121 233 122 234
rect 122 233 123 234
rect 123 233 124 234
rect 124 233 125 234
rect 125 233 126 234
rect 126 233 127 234
rect 127 233 128 234
rect 128 233 129 234
rect 129 233 130 234
rect 130 233 131 234
rect 131 233 132 234
rect 132 233 133 234
rect 133 233 134 234
rect 134 233 135 234
rect 135 233 136 234
rect 136 233 137 234
rect 137 233 138 234
rect 138 233 139 234
rect 139 233 140 234
rect 140 233 141 234
rect 141 233 142 234
rect 142 233 143 234
rect 143 233 144 234
rect 144 233 145 234
rect 145 233 146 234
rect 146 233 147 234
rect 147 233 148 234
rect 148 233 149 234
rect 149 233 150 234
rect 150 233 151 234
rect 151 233 152 234
rect 152 233 153 234
rect 153 233 154 234
rect 154 233 155 234
rect 155 233 156 234
rect 156 233 157 234
rect 157 233 158 234
rect 158 233 159 234
rect 159 233 160 234
rect 160 233 161 234
rect 161 233 162 234
rect 162 233 163 234
rect 163 233 164 234
rect 164 233 165 234
rect 165 233 166 234
rect 166 233 167 234
rect 167 233 168 234
rect 168 233 169 234
rect 169 233 170 234
rect 170 233 171 234
rect 171 233 172 234
rect 172 233 173 234
rect 173 233 174 234
rect 174 233 175 234
rect 186 233 187 234
rect 187 233 188 234
rect 188 233 189 234
rect 189 233 190 234
rect 190 233 191 234
rect 191 233 192 234
rect 192 233 193 234
rect 193 233 194 234
rect 194 233 195 234
rect 195 233 196 234
rect 196 233 197 234
rect 197 233 198 234
rect 198 233 199 234
rect 202 233 203 234
rect 203 233 204 234
rect 204 233 205 234
rect 205 233 206 234
rect 206 233 207 234
rect 207 233 208 234
rect 208 233 209 234
rect 209 233 210 234
rect 210 233 211 234
rect 211 233 212 234
rect 212 233 213 234
rect 213 233 214 234
rect 229 233 230 234
rect 230 233 231 234
rect 231 233 232 234
rect 232 233 233 234
rect 233 233 234 234
rect 234 233 235 234
rect 235 233 236 234
rect 236 233 237 234
rect 237 233 238 234
rect 238 233 239 234
rect 239 233 240 234
rect 240 233 241 234
rect 241 233 242 234
rect 242 233 243 234
rect 243 233 244 234
rect 244 233 245 234
rect 245 233 246 234
rect 246 233 247 234
rect 247 233 248 234
rect 248 233 249 234
rect 249 233 250 234
rect 250 233 251 234
rect 251 233 252 234
rect 252 233 253 234
rect 253 233 254 234
rect 254 233 255 234
rect 255 233 256 234
rect 256 233 257 234
rect 257 233 258 234
rect 258 233 259 234
rect 259 233 260 234
rect 260 233 261 234
rect 261 233 262 234
rect 262 233 263 234
rect 263 233 264 234
rect 264 233 265 234
rect 265 233 266 234
rect 266 233 267 234
rect 267 233 268 234
rect 268 233 269 234
rect 269 233 270 234
rect 270 233 271 234
rect 271 233 272 234
rect 272 233 273 234
rect 273 233 274 234
rect 274 233 275 234
rect 275 233 276 234
rect 276 233 277 234
rect 277 233 278 234
rect 278 233 279 234
rect 279 233 280 234
rect 280 233 281 234
rect 281 233 282 234
rect 282 233 283 234
rect 308 233 309 234
rect 309 233 310 234
rect 310 233 311 234
rect 334 233 335 234
rect 335 233 336 234
rect 336 233 337 234
rect 337 233 338 234
rect 338 233 339 234
rect 363 233 364 234
rect 364 233 365 234
rect 365 233 366 234
rect 366 233 367 234
rect 367 233 368 234
rect 368 233 369 234
rect 369 233 370 234
rect 370 233 371 234
rect 371 233 372 234
rect 372 233 373 234
rect 402 233 403 234
rect 403 233 404 234
rect 404 233 405 234
rect 405 233 406 234
rect 406 233 407 234
rect 407 233 408 234
rect 408 233 409 234
rect 86 232 87 233
rect 87 232 88 233
rect 88 232 89 233
rect 89 232 90 233
rect 90 232 91 233
rect 91 232 92 233
rect 92 232 93 233
rect 93 232 94 233
rect 94 232 95 233
rect 95 232 96 233
rect 96 232 97 233
rect 97 232 98 233
rect 98 232 99 233
rect 99 232 100 233
rect 100 232 101 233
rect 101 232 102 233
rect 102 232 103 233
rect 103 232 104 233
rect 112 232 113 233
rect 113 232 114 233
rect 114 232 115 233
rect 115 232 116 233
rect 116 232 117 233
rect 117 232 118 233
rect 118 232 119 233
rect 119 232 120 233
rect 120 232 121 233
rect 121 232 122 233
rect 122 232 123 233
rect 123 232 124 233
rect 124 232 125 233
rect 125 232 126 233
rect 126 232 127 233
rect 127 232 128 233
rect 128 232 129 233
rect 129 232 130 233
rect 130 232 131 233
rect 131 232 132 233
rect 132 232 133 233
rect 133 232 134 233
rect 134 232 135 233
rect 135 232 136 233
rect 136 232 137 233
rect 137 232 138 233
rect 138 232 139 233
rect 139 232 140 233
rect 140 232 141 233
rect 141 232 142 233
rect 142 232 143 233
rect 143 232 144 233
rect 144 232 145 233
rect 145 232 146 233
rect 146 232 147 233
rect 147 232 148 233
rect 148 232 149 233
rect 149 232 150 233
rect 150 232 151 233
rect 151 232 152 233
rect 152 232 153 233
rect 153 232 154 233
rect 154 232 155 233
rect 155 232 156 233
rect 156 232 157 233
rect 157 232 158 233
rect 158 232 159 233
rect 159 232 160 233
rect 160 232 161 233
rect 161 232 162 233
rect 162 232 163 233
rect 163 232 164 233
rect 164 232 165 233
rect 165 232 166 233
rect 166 232 167 233
rect 167 232 168 233
rect 168 232 169 233
rect 169 232 170 233
rect 170 232 171 233
rect 171 232 172 233
rect 172 232 173 233
rect 173 232 174 233
rect 187 232 188 233
rect 188 232 189 233
rect 189 232 190 233
rect 190 232 191 233
rect 191 232 192 233
rect 192 232 193 233
rect 193 232 194 233
rect 194 232 195 233
rect 195 232 196 233
rect 196 232 197 233
rect 197 232 198 233
rect 198 232 199 233
rect 199 232 200 233
rect 200 232 201 233
rect 201 232 202 233
rect 202 232 203 233
rect 203 232 204 233
rect 204 232 205 233
rect 205 232 206 233
rect 206 232 207 233
rect 207 232 208 233
rect 208 232 209 233
rect 209 232 210 233
rect 210 232 211 233
rect 211 232 212 233
rect 212 232 213 233
rect 230 232 231 233
rect 231 232 232 233
rect 232 232 233 233
rect 233 232 234 233
rect 234 232 235 233
rect 235 232 236 233
rect 236 232 237 233
rect 237 232 238 233
rect 238 232 239 233
rect 239 232 240 233
rect 240 232 241 233
rect 241 232 242 233
rect 242 232 243 233
rect 243 232 244 233
rect 244 232 245 233
rect 245 232 246 233
rect 246 232 247 233
rect 247 232 248 233
rect 248 232 249 233
rect 249 232 250 233
rect 250 232 251 233
rect 251 232 252 233
rect 252 232 253 233
rect 253 232 254 233
rect 254 232 255 233
rect 255 232 256 233
rect 256 232 257 233
rect 257 232 258 233
rect 258 232 259 233
rect 259 232 260 233
rect 260 232 261 233
rect 261 232 262 233
rect 262 232 263 233
rect 263 232 264 233
rect 264 232 265 233
rect 265 232 266 233
rect 266 232 267 233
rect 267 232 268 233
rect 268 232 269 233
rect 269 232 270 233
rect 270 232 271 233
rect 271 232 272 233
rect 272 232 273 233
rect 273 232 274 233
rect 274 232 275 233
rect 275 232 276 233
rect 276 232 277 233
rect 277 232 278 233
rect 278 232 279 233
rect 279 232 280 233
rect 280 232 281 233
rect 281 232 282 233
rect 282 232 283 233
rect 283 232 284 233
rect 284 232 285 233
rect 285 232 286 233
rect 306 232 307 233
rect 307 232 308 233
rect 308 232 309 233
rect 309 232 310 233
rect 334 232 335 233
rect 335 232 336 233
rect 336 232 337 233
rect 337 232 338 233
rect 338 232 339 233
rect 339 232 340 233
rect 361 232 362 233
rect 362 232 363 233
rect 363 232 364 233
rect 364 232 365 233
rect 365 232 366 233
rect 366 232 367 233
rect 367 232 368 233
rect 368 232 369 233
rect 369 232 370 233
rect 370 232 371 233
rect 371 232 372 233
rect 401 232 402 233
rect 402 232 403 233
rect 403 232 404 233
rect 404 232 405 233
rect 405 232 406 233
rect 406 232 407 233
rect 407 232 408 233
rect 87 231 88 232
rect 88 231 89 232
rect 89 231 90 232
rect 90 231 91 232
rect 91 231 92 232
rect 92 231 93 232
rect 93 231 94 232
rect 94 231 95 232
rect 95 231 96 232
rect 96 231 97 232
rect 97 231 98 232
rect 98 231 99 232
rect 99 231 100 232
rect 100 231 101 232
rect 101 231 102 232
rect 102 231 103 232
rect 103 231 104 232
rect 104 231 105 232
rect 105 231 106 232
rect 116 231 117 232
rect 117 231 118 232
rect 118 231 119 232
rect 119 231 120 232
rect 120 231 121 232
rect 121 231 122 232
rect 122 231 123 232
rect 123 231 124 232
rect 124 231 125 232
rect 125 231 126 232
rect 126 231 127 232
rect 127 231 128 232
rect 128 231 129 232
rect 129 231 130 232
rect 130 231 131 232
rect 131 231 132 232
rect 132 231 133 232
rect 133 231 134 232
rect 134 231 135 232
rect 135 231 136 232
rect 136 231 137 232
rect 137 231 138 232
rect 138 231 139 232
rect 139 231 140 232
rect 140 231 141 232
rect 141 231 142 232
rect 142 231 143 232
rect 143 231 144 232
rect 144 231 145 232
rect 145 231 146 232
rect 146 231 147 232
rect 147 231 148 232
rect 148 231 149 232
rect 149 231 150 232
rect 150 231 151 232
rect 151 231 152 232
rect 152 231 153 232
rect 153 231 154 232
rect 154 231 155 232
rect 155 231 156 232
rect 156 231 157 232
rect 157 231 158 232
rect 158 231 159 232
rect 159 231 160 232
rect 160 231 161 232
rect 161 231 162 232
rect 162 231 163 232
rect 163 231 164 232
rect 164 231 165 232
rect 165 231 166 232
rect 166 231 167 232
rect 167 231 168 232
rect 168 231 169 232
rect 169 231 170 232
rect 170 231 171 232
rect 171 231 172 232
rect 172 231 173 232
rect 188 231 189 232
rect 189 231 190 232
rect 190 231 191 232
rect 191 231 192 232
rect 192 231 193 232
rect 193 231 194 232
rect 194 231 195 232
rect 195 231 196 232
rect 196 231 197 232
rect 197 231 198 232
rect 198 231 199 232
rect 199 231 200 232
rect 200 231 201 232
rect 201 231 202 232
rect 202 231 203 232
rect 203 231 204 232
rect 204 231 205 232
rect 205 231 206 232
rect 206 231 207 232
rect 207 231 208 232
rect 208 231 209 232
rect 209 231 210 232
rect 210 231 211 232
rect 211 231 212 232
rect 232 231 233 232
rect 233 231 234 232
rect 234 231 235 232
rect 235 231 236 232
rect 236 231 237 232
rect 237 231 238 232
rect 238 231 239 232
rect 239 231 240 232
rect 240 231 241 232
rect 241 231 242 232
rect 242 231 243 232
rect 243 231 244 232
rect 244 231 245 232
rect 245 231 246 232
rect 246 231 247 232
rect 247 231 248 232
rect 248 231 249 232
rect 249 231 250 232
rect 250 231 251 232
rect 251 231 252 232
rect 252 231 253 232
rect 253 231 254 232
rect 254 231 255 232
rect 255 231 256 232
rect 256 231 257 232
rect 257 231 258 232
rect 258 231 259 232
rect 259 231 260 232
rect 260 231 261 232
rect 261 231 262 232
rect 262 231 263 232
rect 263 231 264 232
rect 264 231 265 232
rect 265 231 266 232
rect 266 231 267 232
rect 267 231 268 232
rect 268 231 269 232
rect 269 231 270 232
rect 270 231 271 232
rect 271 231 272 232
rect 272 231 273 232
rect 273 231 274 232
rect 274 231 275 232
rect 275 231 276 232
rect 276 231 277 232
rect 277 231 278 232
rect 278 231 279 232
rect 279 231 280 232
rect 280 231 281 232
rect 281 231 282 232
rect 282 231 283 232
rect 283 231 284 232
rect 284 231 285 232
rect 285 231 286 232
rect 286 231 287 232
rect 287 231 288 232
rect 288 231 289 232
rect 302 231 303 232
rect 303 231 304 232
rect 304 231 305 232
rect 305 231 306 232
rect 306 231 307 232
rect 307 231 308 232
rect 308 231 309 232
rect 309 231 310 232
rect 334 231 335 232
rect 335 231 336 232
rect 336 231 337 232
rect 337 231 338 232
rect 338 231 339 232
rect 339 231 340 232
rect 340 231 341 232
rect 360 231 361 232
rect 361 231 362 232
rect 362 231 363 232
rect 363 231 364 232
rect 364 231 365 232
rect 365 231 366 232
rect 366 231 367 232
rect 367 231 368 232
rect 368 231 369 232
rect 369 231 370 232
rect 370 231 371 232
rect 401 231 402 232
rect 402 231 403 232
rect 403 231 404 232
rect 404 231 405 232
rect 405 231 406 232
rect 406 231 407 232
rect 407 231 408 232
rect 89 230 90 231
rect 90 230 91 231
rect 91 230 92 231
rect 92 230 93 231
rect 93 230 94 231
rect 94 230 95 231
rect 95 230 96 231
rect 96 230 97 231
rect 97 230 98 231
rect 98 230 99 231
rect 99 230 100 231
rect 100 230 101 231
rect 101 230 102 231
rect 102 230 103 231
rect 103 230 104 231
rect 104 230 105 231
rect 105 230 106 231
rect 106 230 107 231
rect 107 230 108 231
rect 115 230 116 231
rect 116 230 117 231
rect 117 230 118 231
rect 118 230 119 231
rect 119 230 120 231
rect 120 230 121 231
rect 121 230 122 231
rect 122 230 123 231
rect 123 230 124 231
rect 124 230 125 231
rect 125 230 126 231
rect 126 230 127 231
rect 127 230 128 231
rect 128 230 129 231
rect 129 230 130 231
rect 130 230 131 231
rect 131 230 132 231
rect 132 230 133 231
rect 133 230 134 231
rect 134 230 135 231
rect 135 230 136 231
rect 136 230 137 231
rect 137 230 138 231
rect 138 230 139 231
rect 139 230 140 231
rect 140 230 141 231
rect 141 230 142 231
rect 142 230 143 231
rect 143 230 144 231
rect 144 230 145 231
rect 145 230 146 231
rect 146 230 147 231
rect 147 230 148 231
rect 148 230 149 231
rect 149 230 150 231
rect 150 230 151 231
rect 151 230 152 231
rect 152 230 153 231
rect 153 230 154 231
rect 154 230 155 231
rect 155 230 156 231
rect 156 230 157 231
rect 157 230 158 231
rect 158 230 159 231
rect 159 230 160 231
rect 160 230 161 231
rect 161 230 162 231
rect 162 230 163 231
rect 163 230 164 231
rect 164 230 165 231
rect 165 230 166 231
rect 166 230 167 231
rect 167 230 168 231
rect 168 230 169 231
rect 169 230 170 231
rect 170 230 171 231
rect 171 230 172 231
rect 189 230 190 231
rect 190 230 191 231
rect 191 230 192 231
rect 192 230 193 231
rect 193 230 194 231
rect 194 230 195 231
rect 195 230 196 231
rect 196 230 197 231
rect 197 230 198 231
rect 198 230 199 231
rect 199 230 200 231
rect 200 230 201 231
rect 201 230 202 231
rect 202 230 203 231
rect 203 230 204 231
rect 204 230 205 231
rect 205 230 206 231
rect 206 230 207 231
rect 207 230 208 231
rect 208 230 209 231
rect 209 230 210 231
rect 234 230 235 231
rect 235 230 236 231
rect 236 230 237 231
rect 237 230 238 231
rect 238 230 239 231
rect 239 230 240 231
rect 240 230 241 231
rect 241 230 242 231
rect 242 230 243 231
rect 243 230 244 231
rect 244 230 245 231
rect 245 230 246 231
rect 246 230 247 231
rect 247 230 248 231
rect 248 230 249 231
rect 249 230 250 231
rect 250 230 251 231
rect 251 230 252 231
rect 252 230 253 231
rect 253 230 254 231
rect 254 230 255 231
rect 255 230 256 231
rect 256 230 257 231
rect 257 230 258 231
rect 258 230 259 231
rect 259 230 260 231
rect 260 230 261 231
rect 261 230 262 231
rect 262 230 263 231
rect 263 230 264 231
rect 264 230 265 231
rect 265 230 266 231
rect 266 230 267 231
rect 267 230 268 231
rect 268 230 269 231
rect 269 230 270 231
rect 270 230 271 231
rect 271 230 272 231
rect 272 230 273 231
rect 273 230 274 231
rect 274 230 275 231
rect 275 230 276 231
rect 276 230 277 231
rect 277 230 278 231
rect 278 230 279 231
rect 279 230 280 231
rect 280 230 281 231
rect 281 230 282 231
rect 282 230 283 231
rect 283 230 284 231
rect 284 230 285 231
rect 285 230 286 231
rect 286 230 287 231
rect 287 230 288 231
rect 288 230 289 231
rect 289 230 290 231
rect 290 230 291 231
rect 291 230 292 231
rect 292 230 293 231
rect 293 230 294 231
rect 294 230 295 231
rect 295 230 296 231
rect 296 230 297 231
rect 297 230 298 231
rect 298 230 299 231
rect 299 230 300 231
rect 300 230 301 231
rect 301 230 302 231
rect 302 230 303 231
rect 303 230 304 231
rect 304 230 305 231
rect 305 230 306 231
rect 306 230 307 231
rect 307 230 308 231
rect 308 230 309 231
rect 334 230 335 231
rect 335 230 336 231
rect 336 230 337 231
rect 337 230 338 231
rect 338 230 339 231
rect 339 230 340 231
rect 340 230 341 231
rect 341 230 342 231
rect 359 230 360 231
rect 360 230 361 231
rect 361 230 362 231
rect 362 230 363 231
rect 363 230 364 231
rect 364 230 365 231
rect 365 230 366 231
rect 366 230 367 231
rect 367 230 368 231
rect 368 230 369 231
rect 369 230 370 231
rect 400 230 401 231
rect 401 230 402 231
rect 402 230 403 231
rect 403 230 404 231
rect 404 230 405 231
rect 405 230 406 231
rect 406 230 407 231
rect 90 229 91 230
rect 91 229 92 230
rect 92 229 93 230
rect 93 229 94 230
rect 94 229 95 230
rect 95 229 96 230
rect 96 229 97 230
rect 97 229 98 230
rect 98 229 99 230
rect 99 229 100 230
rect 100 229 101 230
rect 101 229 102 230
rect 102 229 103 230
rect 103 229 104 230
rect 104 229 105 230
rect 105 229 106 230
rect 106 229 107 230
rect 107 229 108 230
rect 108 229 109 230
rect 109 229 110 230
rect 110 229 111 230
rect 113 229 114 230
rect 114 229 115 230
rect 115 229 116 230
rect 116 229 117 230
rect 117 229 118 230
rect 118 229 119 230
rect 119 229 120 230
rect 120 229 121 230
rect 121 229 122 230
rect 122 229 123 230
rect 123 229 124 230
rect 124 229 125 230
rect 125 229 126 230
rect 126 229 127 230
rect 127 229 128 230
rect 128 229 129 230
rect 129 229 130 230
rect 130 229 131 230
rect 131 229 132 230
rect 132 229 133 230
rect 133 229 134 230
rect 134 229 135 230
rect 135 229 136 230
rect 136 229 137 230
rect 137 229 138 230
rect 138 229 139 230
rect 139 229 140 230
rect 140 229 141 230
rect 141 229 142 230
rect 142 229 143 230
rect 143 229 144 230
rect 144 229 145 230
rect 145 229 146 230
rect 146 229 147 230
rect 147 229 148 230
rect 148 229 149 230
rect 149 229 150 230
rect 150 229 151 230
rect 151 229 152 230
rect 152 229 153 230
rect 153 229 154 230
rect 154 229 155 230
rect 155 229 156 230
rect 156 229 157 230
rect 157 229 158 230
rect 158 229 159 230
rect 159 229 160 230
rect 160 229 161 230
rect 161 229 162 230
rect 162 229 163 230
rect 163 229 164 230
rect 164 229 165 230
rect 165 229 166 230
rect 166 229 167 230
rect 167 229 168 230
rect 168 229 169 230
rect 169 229 170 230
rect 170 229 171 230
rect 171 229 172 230
rect 191 229 192 230
rect 192 229 193 230
rect 193 229 194 230
rect 194 229 195 230
rect 195 229 196 230
rect 196 229 197 230
rect 197 229 198 230
rect 198 229 199 230
rect 199 229 200 230
rect 200 229 201 230
rect 201 229 202 230
rect 202 229 203 230
rect 203 229 204 230
rect 204 229 205 230
rect 205 229 206 230
rect 206 229 207 230
rect 207 229 208 230
rect 208 229 209 230
rect 235 229 236 230
rect 236 229 237 230
rect 237 229 238 230
rect 238 229 239 230
rect 239 229 240 230
rect 240 229 241 230
rect 241 229 242 230
rect 242 229 243 230
rect 243 229 244 230
rect 244 229 245 230
rect 245 229 246 230
rect 246 229 247 230
rect 247 229 248 230
rect 248 229 249 230
rect 249 229 250 230
rect 250 229 251 230
rect 251 229 252 230
rect 252 229 253 230
rect 253 229 254 230
rect 254 229 255 230
rect 255 229 256 230
rect 256 229 257 230
rect 257 229 258 230
rect 258 229 259 230
rect 259 229 260 230
rect 260 229 261 230
rect 261 229 262 230
rect 262 229 263 230
rect 263 229 264 230
rect 264 229 265 230
rect 265 229 266 230
rect 266 229 267 230
rect 267 229 268 230
rect 268 229 269 230
rect 269 229 270 230
rect 270 229 271 230
rect 271 229 272 230
rect 272 229 273 230
rect 273 229 274 230
rect 274 229 275 230
rect 275 229 276 230
rect 276 229 277 230
rect 277 229 278 230
rect 278 229 279 230
rect 279 229 280 230
rect 280 229 281 230
rect 281 229 282 230
rect 282 229 283 230
rect 283 229 284 230
rect 284 229 285 230
rect 285 229 286 230
rect 286 229 287 230
rect 287 229 288 230
rect 288 229 289 230
rect 289 229 290 230
rect 290 229 291 230
rect 291 229 292 230
rect 292 229 293 230
rect 293 229 294 230
rect 294 229 295 230
rect 295 229 296 230
rect 296 229 297 230
rect 297 229 298 230
rect 298 229 299 230
rect 299 229 300 230
rect 300 229 301 230
rect 301 229 302 230
rect 302 229 303 230
rect 303 229 304 230
rect 304 229 305 230
rect 305 229 306 230
rect 306 229 307 230
rect 307 229 308 230
rect 308 229 309 230
rect 334 229 335 230
rect 335 229 336 230
rect 336 229 337 230
rect 337 229 338 230
rect 338 229 339 230
rect 339 229 340 230
rect 340 229 341 230
rect 341 229 342 230
rect 342 229 343 230
rect 357 229 358 230
rect 358 229 359 230
rect 359 229 360 230
rect 360 229 361 230
rect 361 229 362 230
rect 362 229 363 230
rect 363 229 364 230
rect 364 229 365 230
rect 365 229 366 230
rect 366 229 367 230
rect 367 229 368 230
rect 368 229 369 230
rect 369 229 370 230
rect 370 229 371 230
rect 399 229 400 230
rect 400 229 401 230
rect 401 229 402 230
rect 402 229 403 230
rect 403 229 404 230
rect 404 229 405 230
rect 405 229 406 230
rect 406 229 407 230
rect 92 228 93 229
rect 93 228 94 229
rect 94 228 95 229
rect 95 228 96 229
rect 96 228 97 229
rect 97 228 98 229
rect 98 228 99 229
rect 99 228 100 229
rect 100 228 101 229
rect 101 228 102 229
rect 102 228 103 229
rect 103 228 104 229
rect 104 228 105 229
rect 105 228 106 229
rect 106 228 107 229
rect 107 228 108 229
rect 108 228 109 229
rect 109 228 110 229
rect 110 228 111 229
rect 111 228 112 229
rect 112 228 113 229
rect 113 228 114 229
rect 114 228 115 229
rect 115 228 116 229
rect 116 228 117 229
rect 117 228 118 229
rect 118 228 119 229
rect 119 228 120 229
rect 120 228 121 229
rect 121 228 122 229
rect 122 228 123 229
rect 123 228 124 229
rect 124 228 125 229
rect 125 228 126 229
rect 126 228 127 229
rect 127 228 128 229
rect 128 228 129 229
rect 129 228 130 229
rect 130 228 131 229
rect 131 228 132 229
rect 132 228 133 229
rect 133 228 134 229
rect 134 228 135 229
rect 135 228 136 229
rect 136 228 137 229
rect 137 228 138 229
rect 138 228 139 229
rect 139 228 140 229
rect 140 228 141 229
rect 141 228 142 229
rect 142 228 143 229
rect 143 228 144 229
rect 144 228 145 229
rect 145 228 146 229
rect 146 228 147 229
rect 147 228 148 229
rect 148 228 149 229
rect 149 228 150 229
rect 150 228 151 229
rect 151 228 152 229
rect 152 228 153 229
rect 153 228 154 229
rect 154 228 155 229
rect 155 228 156 229
rect 156 228 157 229
rect 157 228 158 229
rect 158 228 159 229
rect 159 228 160 229
rect 160 228 161 229
rect 161 228 162 229
rect 162 228 163 229
rect 163 228 164 229
rect 164 228 165 229
rect 165 228 166 229
rect 166 228 167 229
rect 167 228 168 229
rect 168 228 169 229
rect 169 228 170 229
rect 170 228 171 229
rect 193 228 194 229
rect 194 228 195 229
rect 195 228 196 229
rect 196 228 197 229
rect 197 228 198 229
rect 198 228 199 229
rect 199 228 200 229
rect 200 228 201 229
rect 201 228 202 229
rect 202 228 203 229
rect 203 228 204 229
rect 204 228 205 229
rect 205 228 206 229
rect 236 228 237 229
rect 237 228 238 229
rect 238 228 239 229
rect 239 228 240 229
rect 240 228 241 229
rect 241 228 242 229
rect 242 228 243 229
rect 243 228 244 229
rect 244 228 245 229
rect 245 228 246 229
rect 246 228 247 229
rect 247 228 248 229
rect 248 228 249 229
rect 249 228 250 229
rect 250 228 251 229
rect 251 228 252 229
rect 252 228 253 229
rect 253 228 254 229
rect 254 228 255 229
rect 255 228 256 229
rect 256 228 257 229
rect 257 228 258 229
rect 258 228 259 229
rect 259 228 260 229
rect 260 228 261 229
rect 261 228 262 229
rect 262 228 263 229
rect 263 228 264 229
rect 264 228 265 229
rect 265 228 266 229
rect 266 228 267 229
rect 267 228 268 229
rect 268 228 269 229
rect 269 228 270 229
rect 270 228 271 229
rect 271 228 272 229
rect 272 228 273 229
rect 273 228 274 229
rect 274 228 275 229
rect 275 228 276 229
rect 276 228 277 229
rect 277 228 278 229
rect 278 228 279 229
rect 279 228 280 229
rect 280 228 281 229
rect 281 228 282 229
rect 282 228 283 229
rect 283 228 284 229
rect 284 228 285 229
rect 285 228 286 229
rect 286 228 287 229
rect 287 228 288 229
rect 288 228 289 229
rect 289 228 290 229
rect 290 228 291 229
rect 291 228 292 229
rect 292 228 293 229
rect 293 228 294 229
rect 294 228 295 229
rect 295 228 296 229
rect 296 228 297 229
rect 297 228 298 229
rect 298 228 299 229
rect 299 228 300 229
rect 300 228 301 229
rect 301 228 302 229
rect 302 228 303 229
rect 303 228 304 229
rect 304 228 305 229
rect 305 228 306 229
rect 306 228 307 229
rect 307 228 308 229
rect 335 228 336 229
rect 336 228 337 229
rect 337 228 338 229
rect 338 228 339 229
rect 339 228 340 229
rect 340 228 341 229
rect 341 228 342 229
rect 342 228 343 229
rect 343 228 344 229
rect 356 228 357 229
rect 357 228 358 229
rect 358 228 359 229
rect 359 228 360 229
rect 360 228 361 229
rect 361 228 362 229
rect 362 228 363 229
rect 363 228 364 229
rect 364 228 365 229
rect 365 228 366 229
rect 366 228 367 229
rect 367 228 368 229
rect 368 228 369 229
rect 369 228 370 229
rect 370 228 371 229
rect 371 228 372 229
rect 372 228 373 229
rect 398 228 399 229
rect 399 228 400 229
rect 400 228 401 229
rect 401 228 402 229
rect 402 228 403 229
rect 403 228 404 229
rect 404 228 405 229
rect 405 228 406 229
rect 94 227 95 228
rect 95 227 96 228
rect 96 227 97 228
rect 97 227 98 228
rect 98 227 99 228
rect 99 227 100 228
rect 100 227 101 228
rect 101 227 102 228
rect 102 227 103 228
rect 103 227 104 228
rect 104 227 105 228
rect 105 227 106 228
rect 106 227 107 228
rect 107 227 108 228
rect 108 227 109 228
rect 109 227 110 228
rect 110 227 111 228
rect 111 227 112 228
rect 112 227 113 228
rect 113 227 114 228
rect 114 227 115 228
rect 115 227 116 228
rect 116 227 117 228
rect 117 227 118 228
rect 118 227 119 228
rect 119 227 120 228
rect 120 227 121 228
rect 121 227 122 228
rect 122 227 123 228
rect 123 227 124 228
rect 124 227 125 228
rect 125 227 126 228
rect 126 227 127 228
rect 127 227 128 228
rect 128 227 129 228
rect 129 227 130 228
rect 130 227 131 228
rect 131 227 132 228
rect 132 227 133 228
rect 133 227 134 228
rect 134 227 135 228
rect 135 227 136 228
rect 136 227 137 228
rect 137 227 138 228
rect 138 227 139 228
rect 139 227 140 228
rect 140 227 141 228
rect 141 227 142 228
rect 142 227 143 228
rect 143 227 144 228
rect 144 227 145 228
rect 145 227 146 228
rect 146 227 147 228
rect 147 227 148 228
rect 148 227 149 228
rect 149 227 150 228
rect 150 227 151 228
rect 151 227 152 228
rect 152 227 153 228
rect 153 227 154 228
rect 154 227 155 228
rect 155 227 156 228
rect 156 227 157 228
rect 157 227 158 228
rect 158 227 159 228
rect 159 227 160 228
rect 160 227 161 228
rect 161 227 162 228
rect 162 227 163 228
rect 163 227 164 228
rect 164 227 165 228
rect 165 227 166 228
rect 166 227 167 228
rect 167 227 168 228
rect 168 227 169 228
rect 169 227 170 228
rect 170 227 171 228
rect 198 227 199 228
rect 199 227 200 228
rect 200 227 201 228
rect 201 227 202 228
rect 238 227 239 228
rect 239 227 240 228
rect 240 227 241 228
rect 241 227 242 228
rect 242 227 243 228
rect 243 227 244 228
rect 244 227 245 228
rect 245 227 246 228
rect 246 227 247 228
rect 247 227 248 228
rect 248 227 249 228
rect 249 227 250 228
rect 250 227 251 228
rect 251 227 252 228
rect 252 227 253 228
rect 253 227 254 228
rect 254 227 255 228
rect 255 227 256 228
rect 256 227 257 228
rect 257 227 258 228
rect 258 227 259 228
rect 259 227 260 228
rect 260 227 261 228
rect 261 227 262 228
rect 262 227 263 228
rect 263 227 264 228
rect 264 227 265 228
rect 265 227 266 228
rect 266 227 267 228
rect 267 227 268 228
rect 268 227 269 228
rect 269 227 270 228
rect 270 227 271 228
rect 271 227 272 228
rect 272 227 273 228
rect 273 227 274 228
rect 274 227 275 228
rect 275 227 276 228
rect 276 227 277 228
rect 277 227 278 228
rect 278 227 279 228
rect 279 227 280 228
rect 280 227 281 228
rect 281 227 282 228
rect 282 227 283 228
rect 283 227 284 228
rect 284 227 285 228
rect 285 227 286 228
rect 286 227 287 228
rect 287 227 288 228
rect 288 227 289 228
rect 289 227 290 228
rect 290 227 291 228
rect 291 227 292 228
rect 292 227 293 228
rect 293 227 294 228
rect 294 227 295 228
rect 295 227 296 228
rect 296 227 297 228
rect 297 227 298 228
rect 298 227 299 228
rect 299 227 300 228
rect 300 227 301 228
rect 301 227 302 228
rect 302 227 303 228
rect 303 227 304 228
rect 304 227 305 228
rect 305 227 306 228
rect 306 227 307 228
rect 335 227 336 228
rect 336 227 337 228
rect 337 227 338 228
rect 338 227 339 228
rect 339 227 340 228
rect 340 227 341 228
rect 341 227 342 228
rect 342 227 343 228
rect 343 227 344 228
rect 344 227 345 228
rect 345 227 346 228
rect 354 227 355 228
rect 355 227 356 228
rect 356 227 357 228
rect 357 227 358 228
rect 358 227 359 228
rect 359 227 360 228
rect 360 227 361 228
rect 361 227 362 228
rect 362 227 363 228
rect 363 227 364 228
rect 364 227 365 228
rect 365 227 366 228
rect 366 227 367 228
rect 367 227 368 228
rect 368 227 369 228
rect 369 227 370 228
rect 370 227 371 228
rect 371 227 372 228
rect 372 227 373 228
rect 373 227 374 228
rect 374 227 375 228
rect 397 227 398 228
rect 398 227 399 228
rect 399 227 400 228
rect 400 227 401 228
rect 401 227 402 228
rect 402 227 403 228
rect 403 227 404 228
rect 404 227 405 228
rect 405 227 406 228
rect 96 226 97 227
rect 97 226 98 227
rect 98 226 99 227
rect 99 226 100 227
rect 100 226 101 227
rect 101 226 102 227
rect 102 226 103 227
rect 103 226 104 227
rect 104 226 105 227
rect 105 226 106 227
rect 106 226 107 227
rect 107 226 108 227
rect 108 226 109 227
rect 109 226 110 227
rect 110 226 111 227
rect 111 226 112 227
rect 112 226 113 227
rect 113 226 114 227
rect 114 226 115 227
rect 115 226 116 227
rect 116 226 117 227
rect 117 226 118 227
rect 118 226 119 227
rect 119 226 120 227
rect 120 226 121 227
rect 121 226 122 227
rect 122 226 123 227
rect 123 226 124 227
rect 124 226 125 227
rect 125 226 126 227
rect 126 226 127 227
rect 127 226 128 227
rect 128 226 129 227
rect 129 226 130 227
rect 130 226 131 227
rect 131 226 132 227
rect 132 226 133 227
rect 133 226 134 227
rect 134 226 135 227
rect 135 226 136 227
rect 136 226 137 227
rect 137 226 138 227
rect 138 226 139 227
rect 139 226 140 227
rect 140 226 141 227
rect 141 226 142 227
rect 142 226 143 227
rect 143 226 144 227
rect 144 226 145 227
rect 145 226 146 227
rect 146 226 147 227
rect 147 226 148 227
rect 148 226 149 227
rect 149 226 150 227
rect 150 226 151 227
rect 151 226 152 227
rect 152 226 153 227
rect 153 226 154 227
rect 154 226 155 227
rect 155 226 156 227
rect 156 226 157 227
rect 157 226 158 227
rect 158 226 159 227
rect 159 226 160 227
rect 160 226 161 227
rect 161 226 162 227
rect 162 226 163 227
rect 163 226 164 227
rect 164 226 165 227
rect 165 226 166 227
rect 166 226 167 227
rect 167 226 168 227
rect 168 226 169 227
rect 169 226 170 227
rect 239 226 240 227
rect 240 226 241 227
rect 241 226 242 227
rect 242 226 243 227
rect 243 226 244 227
rect 244 226 245 227
rect 245 226 246 227
rect 246 226 247 227
rect 247 226 248 227
rect 248 226 249 227
rect 249 226 250 227
rect 250 226 251 227
rect 251 226 252 227
rect 252 226 253 227
rect 253 226 254 227
rect 254 226 255 227
rect 255 226 256 227
rect 256 226 257 227
rect 257 226 258 227
rect 258 226 259 227
rect 259 226 260 227
rect 260 226 261 227
rect 261 226 262 227
rect 262 226 263 227
rect 263 226 264 227
rect 264 226 265 227
rect 265 226 266 227
rect 266 226 267 227
rect 267 226 268 227
rect 268 226 269 227
rect 269 226 270 227
rect 270 226 271 227
rect 271 226 272 227
rect 272 226 273 227
rect 273 226 274 227
rect 274 226 275 227
rect 275 226 276 227
rect 276 226 277 227
rect 277 226 278 227
rect 278 226 279 227
rect 279 226 280 227
rect 280 226 281 227
rect 281 226 282 227
rect 282 226 283 227
rect 283 226 284 227
rect 284 226 285 227
rect 285 226 286 227
rect 286 226 287 227
rect 287 226 288 227
rect 288 226 289 227
rect 289 226 290 227
rect 290 226 291 227
rect 291 226 292 227
rect 292 226 293 227
rect 293 226 294 227
rect 294 226 295 227
rect 295 226 296 227
rect 296 226 297 227
rect 297 226 298 227
rect 298 226 299 227
rect 299 226 300 227
rect 300 226 301 227
rect 301 226 302 227
rect 302 226 303 227
rect 303 226 304 227
rect 304 226 305 227
rect 305 226 306 227
rect 335 226 336 227
rect 336 226 337 227
rect 337 226 338 227
rect 338 226 339 227
rect 339 226 340 227
rect 340 226 341 227
rect 341 226 342 227
rect 342 226 343 227
rect 343 226 344 227
rect 344 226 345 227
rect 345 226 346 227
rect 346 226 347 227
rect 347 226 348 227
rect 348 226 349 227
rect 349 226 350 227
rect 350 226 351 227
rect 351 226 352 227
rect 352 226 353 227
rect 353 226 354 227
rect 354 226 355 227
rect 355 226 356 227
rect 356 226 357 227
rect 357 226 358 227
rect 358 226 359 227
rect 359 226 360 227
rect 360 226 361 227
rect 361 226 362 227
rect 362 226 363 227
rect 363 226 364 227
rect 364 226 365 227
rect 365 226 366 227
rect 366 226 367 227
rect 367 226 368 227
rect 368 226 369 227
rect 369 226 370 227
rect 370 226 371 227
rect 371 226 372 227
rect 372 226 373 227
rect 373 226 374 227
rect 374 226 375 227
rect 375 226 376 227
rect 376 226 377 227
rect 396 226 397 227
rect 397 226 398 227
rect 398 226 399 227
rect 399 226 400 227
rect 400 226 401 227
rect 401 226 402 227
rect 402 226 403 227
rect 403 226 404 227
rect 404 226 405 227
rect 98 225 99 226
rect 99 225 100 226
rect 100 225 101 226
rect 101 225 102 226
rect 102 225 103 226
rect 103 225 104 226
rect 104 225 105 226
rect 105 225 106 226
rect 106 225 107 226
rect 107 225 108 226
rect 108 225 109 226
rect 109 225 110 226
rect 110 225 111 226
rect 111 225 112 226
rect 112 225 113 226
rect 113 225 114 226
rect 114 225 115 226
rect 115 225 116 226
rect 116 225 117 226
rect 117 225 118 226
rect 118 225 119 226
rect 119 225 120 226
rect 120 225 121 226
rect 121 225 122 226
rect 122 225 123 226
rect 123 225 124 226
rect 124 225 125 226
rect 125 225 126 226
rect 126 225 127 226
rect 127 225 128 226
rect 128 225 129 226
rect 129 225 130 226
rect 130 225 131 226
rect 131 225 132 226
rect 132 225 133 226
rect 133 225 134 226
rect 134 225 135 226
rect 135 225 136 226
rect 136 225 137 226
rect 137 225 138 226
rect 138 225 139 226
rect 139 225 140 226
rect 140 225 141 226
rect 141 225 142 226
rect 142 225 143 226
rect 143 225 144 226
rect 144 225 145 226
rect 145 225 146 226
rect 146 225 147 226
rect 147 225 148 226
rect 148 225 149 226
rect 149 225 150 226
rect 150 225 151 226
rect 151 225 152 226
rect 152 225 153 226
rect 153 225 154 226
rect 154 225 155 226
rect 155 225 156 226
rect 156 225 157 226
rect 157 225 158 226
rect 158 225 159 226
rect 159 225 160 226
rect 160 225 161 226
rect 161 225 162 226
rect 162 225 163 226
rect 163 225 164 226
rect 164 225 165 226
rect 165 225 166 226
rect 166 225 167 226
rect 167 225 168 226
rect 168 225 169 226
rect 169 225 170 226
rect 240 225 241 226
rect 241 225 242 226
rect 242 225 243 226
rect 243 225 244 226
rect 244 225 245 226
rect 245 225 246 226
rect 246 225 247 226
rect 247 225 248 226
rect 248 225 249 226
rect 249 225 250 226
rect 250 225 251 226
rect 251 225 252 226
rect 252 225 253 226
rect 253 225 254 226
rect 254 225 255 226
rect 255 225 256 226
rect 256 225 257 226
rect 257 225 258 226
rect 258 225 259 226
rect 259 225 260 226
rect 260 225 261 226
rect 261 225 262 226
rect 262 225 263 226
rect 263 225 264 226
rect 264 225 265 226
rect 265 225 266 226
rect 266 225 267 226
rect 267 225 268 226
rect 268 225 269 226
rect 269 225 270 226
rect 270 225 271 226
rect 271 225 272 226
rect 272 225 273 226
rect 273 225 274 226
rect 274 225 275 226
rect 275 225 276 226
rect 276 225 277 226
rect 277 225 278 226
rect 278 225 279 226
rect 279 225 280 226
rect 280 225 281 226
rect 281 225 282 226
rect 282 225 283 226
rect 283 225 284 226
rect 284 225 285 226
rect 285 225 286 226
rect 286 225 287 226
rect 287 225 288 226
rect 288 225 289 226
rect 289 225 290 226
rect 290 225 291 226
rect 291 225 292 226
rect 292 225 293 226
rect 293 225 294 226
rect 294 225 295 226
rect 295 225 296 226
rect 296 225 297 226
rect 297 225 298 226
rect 298 225 299 226
rect 299 225 300 226
rect 300 225 301 226
rect 301 225 302 226
rect 302 225 303 226
rect 303 225 304 226
rect 304 225 305 226
rect 335 225 336 226
rect 336 225 337 226
rect 337 225 338 226
rect 338 225 339 226
rect 339 225 340 226
rect 340 225 341 226
rect 341 225 342 226
rect 342 225 343 226
rect 343 225 344 226
rect 344 225 345 226
rect 345 225 346 226
rect 346 225 347 226
rect 347 225 348 226
rect 348 225 349 226
rect 349 225 350 226
rect 350 225 351 226
rect 351 225 352 226
rect 352 225 353 226
rect 353 225 354 226
rect 354 225 355 226
rect 355 225 356 226
rect 356 225 357 226
rect 357 225 358 226
rect 358 225 359 226
rect 359 225 360 226
rect 360 225 361 226
rect 361 225 362 226
rect 362 225 363 226
rect 363 225 364 226
rect 364 225 365 226
rect 366 225 367 226
rect 367 225 368 226
rect 368 225 369 226
rect 369 225 370 226
rect 370 225 371 226
rect 371 225 372 226
rect 372 225 373 226
rect 373 225 374 226
rect 374 225 375 226
rect 375 225 376 226
rect 376 225 377 226
rect 377 225 378 226
rect 378 225 379 226
rect 379 225 380 226
rect 394 225 395 226
rect 395 225 396 226
rect 396 225 397 226
rect 397 225 398 226
rect 398 225 399 226
rect 399 225 400 226
rect 400 225 401 226
rect 401 225 402 226
rect 402 225 403 226
rect 403 225 404 226
rect 99 224 100 225
rect 100 224 101 225
rect 101 224 102 225
rect 102 224 103 225
rect 103 224 104 225
rect 104 224 105 225
rect 105 224 106 225
rect 106 224 107 225
rect 107 224 108 225
rect 108 224 109 225
rect 109 224 110 225
rect 110 224 111 225
rect 111 224 112 225
rect 112 224 113 225
rect 113 224 114 225
rect 114 224 115 225
rect 115 224 116 225
rect 116 224 117 225
rect 117 224 118 225
rect 118 224 119 225
rect 119 224 120 225
rect 120 224 121 225
rect 121 224 122 225
rect 122 224 123 225
rect 123 224 124 225
rect 124 224 125 225
rect 125 224 126 225
rect 126 224 127 225
rect 127 224 128 225
rect 128 224 129 225
rect 129 224 130 225
rect 130 224 131 225
rect 131 224 132 225
rect 132 224 133 225
rect 133 224 134 225
rect 134 224 135 225
rect 135 224 136 225
rect 136 224 137 225
rect 137 224 138 225
rect 138 224 139 225
rect 139 224 140 225
rect 140 224 141 225
rect 141 224 142 225
rect 142 224 143 225
rect 143 224 144 225
rect 144 224 145 225
rect 145 224 146 225
rect 146 224 147 225
rect 147 224 148 225
rect 148 224 149 225
rect 149 224 150 225
rect 150 224 151 225
rect 151 224 152 225
rect 152 224 153 225
rect 153 224 154 225
rect 154 224 155 225
rect 155 224 156 225
rect 156 224 157 225
rect 157 224 158 225
rect 158 224 159 225
rect 159 224 160 225
rect 160 224 161 225
rect 163 224 164 225
rect 164 224 165 225
rect 165 224 166 225
rect 166 224 167 225
rect 167 224 168 225
rect 168 224 169 225
rect 241 224 242 225
rect 242 224 243 225
rect 243 224 244 225
rect 244 224 245 225
rect 245 224 246 225
rect 246 224 247 225
rect 247 224 248 225
rect 248 224 249 225
rect 249 224 250 225
rect 250 224 251 225
rect 251 224 252 225
rect 252 224 253 225
rect 253 224 254 225
rect 254 224 255 225
rect 255 224 256 225
rect 256 224 257 225
rect 257 224 258 225
rect 258 224 259 225
rect 259 224 260 225
rect 260 224 261 225
rect 261 224 262 225
rect 262 224 263 225
rect 263 224 264 225
rect 264 224 265 225
rect 265 224 266 225
rect 266 224 267 225
rect 267 224 268 225
rect 268 224 269 225
rect 269 224 270 225
rect 270 224 271 225
rect 271 224 272 225
rect 272 224 273 225
rect 273 224 274 225
rect 274 224 275 225
rect 275 224 276 225
rect 276 224 277 225
rect 277 224 278 225
rect 278 224 279 225
rect 279 224 280 225
rect 280 224 281 225
rect 281 224 282 225
rect 282 224 283 225
rect 283 224 284 225
rect 284 224 285 225
rect 285 224 286 225
rect 286 224 287 225
rect 287 224 288 225
rect 288 224 289 225
rect 289 224 290 225
rect 290 224 291 225
rect 291 224 292 225
rect 292 224 293 225
rect 293 224 294 225
rect 294 224 295 225
rect 295 224 296 225
rect 296 224 297 225
rect 297 224 298 225
rect 298 224 299 225
rect 299 224 300 225
rect 300 224 301 225
rect 301 224 302 225
rect 302 224 303 225
rect 303 224 304 225
rect 335 224 336 225
rect 336 224 337 225
rect 337 224 338 225
rect 338 224 339 225
rect 339 224 340 225
rect 340 224 341 225
rect 341 224 342 225
rect 342 224 343 225
rect 343 224 344 225
rect 344 224 345 225
rect 345 224 346 225
rect 346 224 347 225
rect 347 224 348 225
rect 348 224 349 225
rect 349 224 350 225
rect 350 224 351 225
rect 351 224 352 225
rect 352 224 353 225
rect 353 224 354 225
rect 354 224 355 225
rect 355 224 356 225
rect 356 224 357 225
rect 357 224 358 225
rect 358 224 359 225
rect 359 224 360 225
rect 360 224 361 225
rect 361 224 362 225
rect 362 224 363 225
rect 366 224 367 225
rect 367 224 368 225
rect 368 224 369 225
rect 369 224 370 225
rect 370 224 371 225
rect 371 224 372 225
rect 372 224 373 225
rect 373 224 374 225
rect 374 224 375 225
rect 375 224 376 225
rect 376 224 377 225
rect 377 224 378 225
rect 378 224 379 225
rect 379 224 380 225
rect 380 224 381 225
rect 381 224 382 225
rect 382 224 383 225
rect 383 224 384 225
rect 391 224 392 225
rect 392 224 393 225
rect 393 224 394 225
rect 394 224 395 225
rect 395 224 396 225
rect 396 224 397 225
rect 397 224 398 225
rect 398 224 399 225
rect 399 224 400 225
rect 400 224 401 225
rect 401 224 402 225
rect 402 224 403 225
rect 403 224 404 225
rect 96 223 97 224
rect 97 223 98 224
rect 98 223 99 224
rect 99 223 100 224
rect 100 223 101 224
rect 101 223 102 224
rect 102 223 103 224
rect 103 223 104 224
rect 104 223 105 224
rect 105 223 106 224
rect 106 223 107 224
rect 107 223 108 224
rect 108 223 109 224
rect 109 223 110 224
rect 110 223 111 224
rect 111 223 112 224
rect 112 223 113 224
rect 113 223 114 224
rect 114 223 115 224
rect 115 223 116 224
rect 116 223 117 224
rect 117 223 118 224
rect 118 223 119 224
rect 119 223 120 224
rect 120 223 121 224
rect 121 223 122 224
rect 122 223 123 224
rect 123 223 124 224
rect 124 223 125 224
rect 125 223 126 224
rect 126 223 127 224
rect 127 223 128 224
rect 128 223 129 224
rect 129 223 130 224
rect 130 223 131 224
rect 131 223 132 224
rect 132 223 133 224
rect 133 223 134 224
rect 134 223 135 224
rect 135 223 136 224
rect 136 223 137 224
rect 137 223 138 224
rect 138 223 139 224
rect 139 223 140 224
rect 140 223 141 224
rect 141 223 142 224
rect 142 223 143 224
rect 143 223 144 224
rect 144 223 145 224
rect 145 223 146 224
rect 146 223 147 224
rect 147 223 148 224
rect 148 223 149 224
rect 149 223 150 224
rect 150 223 151 224
rect 151 223 152 224
rect 152 223 153 224
rect 153 223 154 224
rect 154 223 155 224
rect 155 223 156 224
rect 156 223 157 224
rect 157 223 158 224
rect 158 223 159 224
rect 159 223 160 224
rect 163 223 164 224
rect 164 223 165 224
rect 165 223 166 224
rect 166 223 167 224
rect 167 223 168 224
rect 168 223 169 224
rect 242 223 243 224
rect 243 223 244 224
rect 244 223 245 224
rect 245 223 246 224
rect 246 223 247 224
rect 247 223 248 224
rect 248 223 249 224
rect 249 223 250 224
rect 250 223 251 224
rect 251 223 252 224
rect 252 223 253 224
rect 253 223 254 224
rect 254 223 255 224
rect 255 223 256 224
rect 256 223 257 224
rect 257 223 258 224
rect 258 223 259 224
rect 259 223 260 224
rect 260 223 261 224
rect 261 223 262 224
rect 262 223 263 224
rect 263 223 264 224
rect 264 223 265 224
rect 265 223 266 224
rect 266 223 267 224
rect 267 223 268 224
rect 268 223 269 224
rect 269 223 270 224
rect 270 223 271 224
rect 271 223 272 224
rect 272 223 273 224
rect 273 223 274 224
rect 274 223 275 224
rect 275 223 276 224
rect 276 223 277 224
rect 277 223 278 224
rect 278 223 279 224
rect 279 223 280 224
rect 280 223 281 224
rect 281 223 282 224
rect 282 223 283 224
rect 283 223 284 224
rect 284 223 285 224
rect 285 223 286 224
rect 286 223 287 224
rect 287 223 288 224
rect 288 223 289 224
rect 289 223 290 224
rect 290 223 291 224
rect 291 223 292 224
rect 292 223 293 224
rect 293 223 294 224
rect 294 223 295 224
rect 295 223 296 224
rect 296 223 297 224
rect 297 223 298 224
rect 298 223 299 224
rect 299 223 300 224
rect 300 223 301 224
rect 301 223 302 224
rect 335 223 336 224
rect 336 223 337 224
rect 337 223 338 224
rect 338 223 339 224
rect 339 223 340 224
rect 340 223 341 224
rect 341 223 342 224
rect 342 223 343 224
rect 343 223 344 224
rect 344 223 345 224
rect 345 223 346 224
rect 346 223 347 224
rect 347 223 348 224
rect 348 223 349 224
rect 349 223 350 224
rect 350 223 351 224
rect 351 223 352 224
rect 352 223 353 224
rect 353 223 354 224
rect 354 223 355 224
rect 355 223 356 224
rect 356 223 357 224
rect 357 223 358 224
rect 358 223 359 224
rect 359 223 360 224
rect 360 223 361 224
rect 361 223 362 224
rect 366 223 367 224
rect 367 223 368 224
rect 368 223 369 224
rect 369 223 370 224
rect 370 223 371 224
rect 371 223 372 224
rect 372 223 373 224
rect 373 223 374 224
rect 374 223 375 224
rect 375 223 376 224
rect 376 223 377 224
rect 377 223 378 224
rect 378 223 379 224
rect 379 223 380 224
rect 380 223 381 224
rect 381 223 382 224
rect 382 223 383 224
rect 383 223 384 224
rect 384 223 385 224
rect 385 223 386 224
rect 386 223 387 224
rect 387 223 388 224
rect 388 223 389 224
rect 389 223 390 224
rect 390 223 391 224
rect 391 223 392 224
rect 392 223 393 224
rect 393 223 394 224
rect 394 223 395 224
rect 395 223 396 224
rect 396 223 397 224
rect 397 223 398 224
rect 398 223 399 224
rect 399 223 400 224
rect 400 223 401 224
rect 401 223 402 224
rect 402 223 403 224
rect 100 222 101 223
rect 101 222 102 223
rect 102 222 103 223
rect 103 222 104 223
rect 104 222 105 223
rect 105 222 106 223
rect 106 222 107 223
rect 107 222 108 223
rect 108 222 109 223
rect 109 222 110 223
rect 110 222 111 223
rect 111 222 112 223
rect 112 222 113 223
rect 113 222 114 223
rect 114 222 115 223
rect 115 222 116 223
rect 116 222 117 223
rect 117 222 118 223
rect 118 222 119 223
rect 119 222 120 223
rect 120 222 121 223
rect 121 222 122 223
rect 122 222 123 223
rect 123 222 124 223
rect 124 222 125 223
rect 125 222 126 223
rect 126 222 127 223
rect 127 222 128 223
rect 128 222 129 223
rect 129 222 130 223
rect 130 222 131 223
rect 131 222 132 223
rect 132 222 133 223
rect 133 222 134 223
rect 134 222 135 223
rect 135 222 136 223
rect 136 222 137 223
rect 137 222 138 223
rect 138 222 139 223
rect 139 222 140 223
rect 140 222 141 223
rect 141 222 142 223
rect 142 222 143 223
rect 143 222 144 223
rect 144 222 145 223
rect 145 222 146 223
rect 146 222 147 223
rect 147 222 148 223
rect 148 222 149 223
rect 149 222 150 223
rect 150 222 151 223
rect 151 222 152 223
rect 152 222 153 223
rect 153 222 154 223
rect 154 222 155 223
rect 155 222 156 223
rect 156 222 157 223
rect 157 222 158 223
rect 163 222 164 223
rect 164 222 165 223
rect 165 222 166 223
rect 166 222 167 223
rect 167 222 168 223
rect 168 222 169 223
rect 243 222 244 223
rect 244 222 245 223
rect 245 222 246 223
rect 246 222 247 223
rect 247 222 248 223
rect 248 222 249 223
rect 249 222 250 223
rect 250 222 251 223
rect 251 222 252 223
rect 252 222 253 223
rect 253 222 254 223
rect 254 222 255 223
rect 255 222 256 223
rect 256 222 257 223
rect 257 222 258 223
rect 258 222 259 223
rect 259 222 260 223
rect 260 222 261 223
rect 261 222 262 223
rect 262 222 263 223
rect 263 222 264 223
rect 264 222 265 223
rect 265 222 266 223
rect 266 222 267 223
rect 267 222 268 223
rect 268 222 269 223
rect 269 222 270 223
rect 270 222 271 223
rect 271 222 272 223
rect 272 222 273 223
rect 273 222 274 223
rect 274 222 275 223
rect 275 222 276 223
rect 276 222 277 223
rect 277 222 278 223
rect 278 222 279 223
rect 279 222 280 223
rect 280 222 281 223
rect 281 222 282 223
rect 282 222 283 223
rect 283 222 284 223
rect 284 222 285 223
rect 285 222 286 223
rect 286 222 287 223
rect 287 222 288 223
rect 288 222 289 223
rect 289 222 290 223
rect 290 222 291 223
rect 291 222 292 223
rect 292 222 293 223
rect 293 222 294 223
rect 294 222 295 223
rect 295 222 296 223
rect 296 222 297 223
rect 297 222 298 223
rect 298 222 299 223
rect 299 222 300 223
rect 335 222 336 223
rect 336 222 337 223
rect 337 222 338 223
rect 338 222 339 223
rect 339 222 340 223
rect 340 222 341 223
rect 341 222 342 223
rect 342 222 343 223
rect 343 222 344 223
rect 344 222 345 223
rect 345 222 346 223
rect 346 222 347 223
rect 347 222 348 223
rect 348 222 349 223
rect 349 222 350 223
rect 350 222 351 223
rect 351 222 352 223
rect 352 222 353 223
rect 353 222 354 223
rect 354 222 355 223
rect 355 222 356 223
rect 356 222 357 223
rect 357 222 358 223
rect 358 222 359 223
rect 359 222 360 223
rect 360 222 361 223
rect 366 222 367 223
rect 367 222 368 223
rect 368 222 369 223
rect 369 222 370 223
rect 370 222 371 223
rect 371 222 372 223
rect 372 222 373 223
rect 373 222 374 223
rect 374 222 375 223
rect 375 222 376 223
rect 376 222 377 223
rect 377 222 378 223
rect 378 222 379 223
rect 379 222 380 223
rect 380 222 381 223
rect 381 222 382 223
rect 382 222 383 223
rect 383 222 384 223
rect 384 222 385 223
rect 385 222 386 223
rect 386 222 387 223
rect 387 222 388 223
rect 388 222 389 223
rect 389 222 390 223
rect 390 222 391 223
rect 391 222 392 223
rect 392 222 393 223
rect 393 222 394 223
rect 394 222 395 223
rect 395 222 396 223
rect 396 222 397 223
rect 397 222 398 223
rect 398 222 399 223
rect 399 222 400 223
rect 400 222 401 223
rect 401 222 402 223
rect 106 221 107 222
rect 107 221 108 222
rect 108 221 109 222
rect 109 221 110 222
rect 110 221 111 222
rect 111 221 112 222
rect 112 221 113 222
rect 113 221 114 222
rect 114 221 115 222
rect 115 221 116 222
rect 116 221 117 222
rect 117 221 118 222
rect 118 221 119 222
rect 119 221 120 222
rect 120 221 121 222
rect 121 221 122 222
rect 122 221 123 222
rect 123 221 124 222
rect 124 221 125 222
rect 125 221 126 222
rect 126 221 127 222
rect 127 221 128 222
rect 128 221 129 222
rect 129 221 130 222
rect 130 221 131 222
rect 131 221 132 222
rect 132 221 133 222
rect 133 221 134 222
rect 134 221 135 222
rect 135 221 136 222
rect 136 221 137 222
rect 137 221 138 222
rect 138 221 139 222
rect 139 221 140 222
rect 140 221 141 222
rect 141 221 142 222
rect 142 221 143 222
rect 143 221 144 222
rect 144 221 145 222
rect 145 221 146 222
rect 146 221 147 222
rect 147 221 148 222
rect 148 221 149 222
rect 149 221 150 222
rect 150 221 151 222
rect 151 221 152 222
rect 152 221 153 222
rect 153 221 154 222
rect 154 221 155 222
rect 155 221 156 222
rect 156 221 157 222
rect 163 221 164 222
rect 164 221 165 222
rect 165 221 166 222
rect 166 221 167 222
rect 167 221 168 222
rect 244 221 245 222
rect 245 221 246 222
rect 246 221 247 222
rect 247 221 248 222
rect 248 221 249 222
rect 249 221 250 222
rect 250 221 251 222
rect 251 221 252 222
rect 252 221 253 222
rect 253 221 254 222
rect 254 221 255 222
rect 255 221 256 222
rect 256 221 257 222
rect 257 221 258 222
rect 258 221 259 222
rect 259 221 260 222
rect 260 221 261 222
rect 261 221 262 222
rect 262 221 263 222
rect 263 221 264 222
rect 264 221 265 222
rect 265 221 266 222
rect 266 221 267 222
rect 267 221 268 222
rect 268 221 269 222
rect 269 221 270 222
rect 270 221 271 222
rect 271 221 272 222
rect 272 221 273 222
rect 273 221 274 222
rect 274 221 275 222
rect 275 221 276 222
rect 276 221 277 222
rect 277 221 278 222
rect 278 221 279 222
rect 279 221 280 222
rect 280 221 281 222
rect 281 221 282 222
rect 282 221 283 222
rect 283 221 284 222
rect 284 221 285 222
rect 285 221 286 222
rect 286 221 287 222
rect 287 221 288 222
rect 288 221 289 222
rect 289 221 290 222
rect 290 221 291 222
rect 291 221 292 222
rect 292 221 293 222
rect 293 221 294 222
rect 294 221 295 222
rect 295 221 296 222
rect 296 221 297 222
rect 297 221 298 222
rect 335 221 336 222
rect 336 221 337 222
rect 337 221 338 222
rect 338 221 339 222
rect 339 221 340 222
rect 341 221 342 222
rect 342 221 343 222
rect 343 221 344 222
rect 344 221 345 222
rect 345 221 346 222
rect 346 221 347 222
rect 347 221 348 222
rect 348 221 349 222
rect 349 221 350 222
rect 350 221 351 222
rect 351 221 352 222
rect 352 221 353 222
rect 353 221 354 222
rect 354 221 355 222
rect 355 221 356 222
rect 356 221 357 222
rect 357 221 358 222
rect 358 221 359 222
rect 359 221 360 222
rect 360 221 361 222
rect 361 221 362 222
rect 366 221 367 222
rect 367 221 368 222
rect 368 221 369 222
rect 369 221 370 222
rect 370 221 371 222
rect 372 221 373 222
rect 373 221 374 222
rect 374 221 375 222
rect 375 221 376 222
rect 376 221 377 222
rect 377 221 378 222
rect 378 221 379 222
rect 379 221 380 222
rect 380 221 381 222
rect 381 221 382 222
rect 382 221 383 222
rect 383 221 384 222
rect 384 221 385 222
rect 385 221 386 222
rect 386 221 387 222
rect 387 221 388 222
rect 388 221 389 222
rect 389 221 390 222
rect 390 221 391 222
rect 391 221 392 222
rect 392 221 393 222
rect 393 221 394 222
rect 394 221 395 222
rect 395 221 396 222
rect 396 221 397 222
rect 397 221 398 222
rect 398 221 399 222
rect 399 221 400 222
rect 111 220 112 221
rect 112 220 113 221
rect 113 220 114 221
rect 114 220 115 221
rect 115 220 116 221
rect 116 220 117 221
rect 117 220 118 221
rect 118 220 119 221
rect 119 220 120 221
rect 120 220 121 221
rect 121 220 122 221
rect 122 220 123 221
rect 123 220 124 221
rect 124 220 125 221
rect 125 220 126 221
rect 126 220 127 221
rect 127 220 128 221
rect 128 220 129 221
rect 129 220 130 221
rect 130 220 131 221
rect 131 220 132 221
rect 132 220 133 221
rect 133 220 134 221
rect 134 220 135 221
rect 135 220 136 221
rect 136 220 137 221
rect 137 220 138 221
rect 138 220 139 221
rect 139 220 140 221
rect 140 220 141 221
rect 141 220 142 221
rect 142 220 143 221
rect 143 220 144 221
rect 144 220 145 221
rect 145 220 146 221
rect 146 220 147 221
rect 147 220 148 221
rect 148 220 149 221
rect 149 220 150 221
rect 150 220 151 221
rect 151 220 152 221
rect 152 220 153 221
rect 153 220 154 221
rect 154 220 155 221
rect 163 220 164 221
rect 164 220 165 221
rect 165 220 166 221
rect 166 220 167 221
rect 167 220 168 221
rect 245 220 246 221
rect 246 220 247 221
rect 247 220 248 221
rect 248 220 249 221
rect 249 220 250 221
rect 250 220 251 221
rect 251 220 252 221
rect 252 220 253 221
rect 253 220 254 221
rect 254 220 255 221
rect 255 220 256 221
rect 256 220 257 221
rect 257 220 258 221
rect 258 220 259 221
rect 259 220 260 221
rect 260 220 261 221
rect 261 220 262 221
rect 262 220 263 221
rect 263 220 264 221
rect 264 220 265 221
rect 265 220 266 221
rect 266 220 267 221
rect 267 220 268 221
rect 268 220 269 221
rect 269 220 270 221
rect 270 220 271 221
rect 271 220 272 221
rect 272 220 273 221
rect 273 220 274 221
rect 274 220 275 221
rect 275 220 276 221
rect 276 220 277 221
rect 277 220 278 221
rect 278 220 279 221
rect 279 220 280 221
rect 280 220 281 221
rect 281 220 282 221
rect 282 220 283 221
rect 283 220 284 221
rect 284 220 285 221
rect 285 220 286 221
rect 286 220 287 221
rect 287 220 288 221
rect 288 220 289 221
rect 289 220 290 221
rect 290 220 291 221
rect 291 220 292 221
rect 292 220 293 221
rect 293 220 294 221
rect 294 220 295 221
rect 335 220 336 221
rect 336 220 337 221
rect 337 220 338 221
rect 338 220 339 221
rect 339 220 340 221
rect 343 220 344 221
rect 344 220 345 221
rect 345 220 346 221
rect 346 220 347 221
rect 347 220 348 221
rect 348 220 349 221
rect 349 220 350 221
rect 350 220 351 221
rect 351 220 352 221
rect 352 220 353 221
rect 353 220 354 221
rect 354 220 355 221
rect 355 220 356 221
rect 356 220 357 221
rect 359 220 360 221
rect 360 220 361 221
rect 361 220 362 221
rect 362 220 363 221
rect 366 220 367 221
rect 367 220 368 221
rect 368 220 369 221
rect 369 220 370 221
rect 370 220 371 221
rect 375 220 376 221
rect 376 220 377 221
rect 377 220 378 221
rect 378 220 379 221
rect 379 220 380 221
rect 380 220 381 221
rect 381 220 382 221
rect 382 220 383 221
rect 383 220 384 221
rect 384 220 385 221
rect 385 220 386 221
rect 386 220 387 221
rect 387 220 388 221
rect 388 220 389 221
rect 389 220 390 221
rect 390 220 391 221
rect 391 220 392 221
rect 392 220 393 221
rect 393 220 394 221
rect 394 220 395 221
rect 395 220 396 221
rect 396 220 397 221
rect 397 220 398 221
rect 398 220 399 221
rect 110 219 111 220
rect 111 219 112 220
rect 112 219 113 220
rect 113 219 114 220
rect 114 219 115 220
rect 115 219 116 220
rect 116 219 117 220
rect 117 219 118 220
rect 118 219 119 220
rect 119 219 120 220
rect 120 219 121 220
rect 121 219 122 220
rect 122 219 123 220
rect 123 219 124 220
rect 124 219 125 220
rect 125 219 126 220
rect 126 219 127 220
rect 127 219 128 220
rect 128 219 129 220
rect 129 219 130 220
rect 130 219 131 220
rect 131 219 132 220
rect 132 219 133 220
rect 133 219 134 220
rect 134 219 135 220
rect 135 219 136 220
rect 136 219 137 220
rect 137 219 138 220
rect 138 219 139 220
rect 139 219 140 220
rect 140 219 141 220
rect 141 219 142 220
rect 142 219 143 220
rect 143 219 144 220
rect 144 219 145 220
rect 145 219 146 220
rect 146 219 147 220
rect 147 219 148 220
rect 148 219 149 220
rect 149 219 150 220
rect 150 219 151 220
rect 151 219 152 220
rect 152 219 153 220
rect 163 219 164 220
rect 164 219 165 220
rect 165 219 166 220
rect 166 219 167 220
rect 167 219 168 220
rect 246 219 247 220
rect 247 219 248 220
rect 248 219 249 220
rect 249 219 250 220
rect 250 219 251 220
rect 251 219 252 220
rect 252 219 253 220
rect 253 219 254 220
rect 254 219 255 220
rect 255 219 256 220
rect 256 219 257 220
rect 257 219 258 220
rect 258 219 259 220
rect 259 219 260 220
rect 260 219 261 220
rect 261 219 262 220
rect 262 219 263 220
rect 263 219 264 220
rect 264 219 265 220
rect 265 219 266 220
rect 266 219 267 220
rect 267 219 268 220
rect 268 219 269 220
rect 269 219 270 220
rect 270 219 271 220
rect 271 219 272 220
rect 272 219 273 220
rect 273 219 274 220
rect 274 219 275 220
rect 275 219 276 220
rect 276 219 277 220
rect 277 219 278 220
rect 278 219 279 220
rect 279 219 280 220
rect 280 219 281 220
rect 281 219 282 220
rect 282 219 283 220
rect 283 219 284 220
rect 284 219 285 220
rect 285 219 286 220
rect 286 219 287 220
rect 287 219 288 220
rect 288 219 289 220
rect 289 219 290 220
rect 290 219 291 220
rect 335 219 336 220
rect 336 219 337 220
rect 337 219 338 220
rect 338 219 339 220
rect 339 219 340 220
rect 346 219 347 220
rect 347 219 348 220
rect 348 219 349 220
rect 349 219 350 220
rect 350 219 351 220
rect 351 219 352 220
rect 352 219 353 220
rect 353 219 354 220
rect 359 219 360 220
rect 360 219 361 220
rect 361 219 362 220
rect 362 219 363 220
rect 363 219 364 220
rect 365 219 366 220
rect 366 219 367 220
rect 367 219 368 220
rect 368 219 369 220
rect 369 219 370 220
rect 377 219 378 220
rect 378 219 379 220
rect 379 219 380 220
rect 380 219 381 220
rect 381 219 382 220
rect 382 219 383 220
rect 383 219 384 220
rect 384 219 385 220
rect 385 219 386 220
rect 386 219 387 220
rect 387 219 388 220
rect 388 219 389 220
rect 389 219 390 220
rect 390 219 391 220
rect 391 219 392 220
rect 392 219 393 220
rect 393 219 394 220
rect 394 219 395 220
rect 395 219 396 220
rect 396 219 397 220
rect 104 218 105 219
rect 105 218 106 219
rect 106 218 107 219
rect 107 218 108 219
rect 108 218 109 219
rect 109 218 110 219
rect 110 218 111 219
rect 111 218 112 219
rect 112 218 113 219
rect 113 218 114 219
rect 114 218 115 219
rect 115 218 116 219
rect 116 218 117 219
rect 117 218 118 219
rect 118 218 119 219
rect 119 218 120 219
rect 120 218 121 219
rect 121 218 122 219
rect 122 218 123 219
rect 123 218 124 219
rect 124 218 125 219
rect 125 218 126 219
rect 126 218 127 219
rect 127 218 128 219
rect 128 218 129 219
rect 129 218 130 219
rect 130 218 131 219
rect 131 218 132 219
rect 132 218 133 219
rect 133 218 134 219
rect 134 218 135 219
rect 135 218 136 219
rect 136 218 137 219
rect 137 218 138 219
rect 138 218 139 219
rect 139 218 140 219
rect 140 218 141 219
rect 141 218 142 219
rect 142 218 143 219
rect 143 218 144 219
rect 144 218 145 219
rect 145 218 146 219
rect 146 218 147 219
rect 147 218 148 219
rect 148 218 149 219
rect 149 218 150 219
rect 163 218 164 219
rect 164 218 165 219
rect 165 218 166 219
rect 166 218 167 219
rect 167 218 168 219
rect 247 218 248 219
rect 248 218 249 219
rect 249 218 250 219
rect 250 218 251 219
rect 251 218 252 219
rect 252 218 253 219
rect 253 218 254 219
rect 254 218 255 219
rect 255 218 256 219
rect 256 218 257 219
rect 257 218 258 219
rect 258 218 259 219
rect 259 218 260 219
rect 260 218 261 219
rect 261 218 262 219
rect 262 218 263 219
rect 263 218 264 219
rect 264 218 265 219
rect 265 218 266 219
rect 266 218 267 219
rect 267 218 268 219
rect 268 218 269 219
rect 269 218 270 219
rect 270 218 271 219
rect 271 218 272 219
rect 272 218 273 219
rect 273 218 274 219
rect 274 218 275 219
rect 275 218 276 219
rect 276 218 277 219
rect 277 218 278 219
rect 278 218 279 219
rect 279 218 280 219
rect 280 218 281 219
rect 281 218 282 219
rect 282 218 283 219
rect 283 218 284 219
rect 284 218 285 219
rect 285 218 286 219
rect 286 218 287 219
rect 287 218 288 219
rect 335 218 336 219
rect 336 218 337 219
rect 337 218 338 219
rect 338 218 339 219
rect 339 218 340 219
rect 360 218 361 219
rect 361 218 362 219
rect 362 218 363 219
rect 363 218 364 219
rect 364 218 365 219
rect 365 218 366 219
rect 366 218 367 219
rect 367 218 368 219
rect 368 218 369 219
rect 369 218 370 219
rect 380 218 381 219
rect 381 218 382 219
rect 382 218 383 219
rect 383 218 384 219
rect 384 218 385 219
rect 385 218 386 219
rect 386 218 387 219
rect 387 218 388 219
rect 388 218 389 219
rect 389 218 390 219
rect 390 218 391 219
rect 391 218 392 219
rect 392 218 393 219
rect 393 218 394 219
rect 96 217 97 218
rect 97 217 98 218
rect 98 217 99 218
rect 99 217 100 218
rect 100 217 101 218
rect 101 217 102 218
rect 102 217 103 218
rect 103 217 104 218
rect 104 217 105 218
rect 105 217 106 218
rect 106 217 107 218
rect 107 217 108 218
rect 108 217 109 218
rect 109 217 110 218
rect 110 217 111 218
rect 111 217 112 218
rect 112 217 113 218
rect 113 217 114 218
rect 114 217 115 218
rect 115 217 116 218
rect 116 217 117 218
rect 117 217 118 218
rect 118 217 119 218
rect 119 217 120 218
rect 120 217 121 218
rect 121 217 122 218
rect 122 217 123 218
rect 123 217 124 218
rect 124 217 125 218
rect 125 217 126 218
rect 126 217 127 218
rect 127 217 128 218
rect 128 217 129 218
rect 129 217 130 218
rect 130 217 131 218
rect 131 217 132 218
rect 132 217 133 218
rect 133 217 134 218
rect 134 217 135 218
rect 135 217 136 218
rect 136 217 137 218
rect 137 217 138 218
rect 138 217 139 218
rect 139 217 140 218
rect 140 217 141 218
rect 141 217 142 218
rect 142 217 143 218
rect 143 217 144 218
rect 144 217 145 218
rect 145 217 146 218
rect 146 217 147 218
rect 147 217 148 218
rect 163 217 164 218
rect 164 217 165 218
rect 165 217 166 218
rect 166 217 167 218
rect 248 217 249 218
rect 249 217 250 218
rect 250 217 251 218
rect 251 217 252 218
rect 252 217 253 218
rect 253 217 254 218
rect 254 217 255 218
rect 255 217 256 218
rect 256 217 257 218
rect 257 217 258 218
rect 258 217 259 218
rect 259 217 260 218
rect 260 217 261 218
rect 261 217 262 218
rect 262 217 263 218
rect 263 217 264 218
rect 264 217 265 218
rect 265 217 266 218
rect 266 217 267 218
rect 267 217 268 218
rect 268 217 269 218
rect 269 217 270 218
rect 270 217 271 218
rect 271 217 272 218
rect 272 217 273 218
rect 273 217 274 218
rect 274 217 275 218
rect 275 217 276 218
rect 276 217 277 218
rect 277 217 278 218
rect 278 217 279 218
rect 279 217 280 218
rect 280 217 281 218
rect 281 217 282 218
rect 282 217 283 218
rect 283 217 284 218
rect 284 217 285 218
rect 285 217 286 218
rect 286 217 287 218
rect 287 217 288 218
rect 335 217 336 218
rect 336 217 337 218
rect 337 217 338 218
rect 338 217 339 218
rect 339 217 340 218
rect 361 217 362 218
rect 362 217 363 218
rect 363 217 364 218
rect 364 217 365 218
rect 365 217 366 218
rect 366 217 367 218
rect 367 217 368 218
rect 368 217 369 218
rect 386 217 387 218
rect 387 217 388 218
rect 388 217 389 218
rect 389 217 390 218
rect 101 216 102 217
rect 102 216 103 217
rect 103 216 104 217
rect 104 216 105 217
rect 105 216 106 217
rect 106 216 107 217
rect 107 216 108 217
rect 108 216 109 217
rect 109 216 110 217
rect 110 216 111 217
rect 111 216 112 217
rect 112 216 113 217
rect 113 216 114 217
rect 114 216 115 217
rect 115 216 116 217
rect 116 216 117 217
rect 117 216 118 217
rect 118 216 119 217
rect 119 216 120 217
rect 120 216 121 217
rect 121 216 122 217
rect 122 216 123 217
rect 123 216 124 217
rect 124 216 125 217
rect 125 216 126 217
rect 126 216 127 217
rect 127 216 128 217
rect 128 216 129 217
rect 129 216 130 217
rect 130 216 131 217
rect 131 216 132 217
rect 132 216 133 217
rect 133 216 134 217
rect 134 216 135 217
rect 135 216 136 217
rect 136 216 137 217
rect 137 216 138 217
rect 138 216 139 217
rect 139 216 140 217
rect 140 216 141 217
rect 141 216 142 217
rect 142 216 143 217
rect 143 216 144 217
rect 144 216 145 217
rect 145 216 146 217
rect 146 216 147 217
rect 163 216 164 217
rect 164 216 165 217
rect 165 216 166 217
rect 166 216 167 217
rect 184 216 185 217
rect 185 216 186 217
rect 186 216 187 217
rect 187 216 188 217
rect 188 216 189 217
rect 189 216 190 217
rect 190 216 191 217
rect 191 216 192 217
rect 192 216 193 217
rect 193 216 194 217
rect 194 216 195 217
rect 249 216 250 217
rect 250 216 251 217
rect 251 216 252 217
rect 252 216 253 217
rect 253 216 254 217
rect 254 216 255 217
rect 255 216 256 217
rect 256 216 257 217
rect 257 216 258 217
rect 258 216 259 217
rect 259 216 260 217
rect 260 216 261 217
rect 261 216 262 217
rect 262 216 263 217
rect 263 216 264 217
rect 264 216 265 217
rect 265 216 266 217
rect 266 216 267 217
rect 267 216 268 217
rect 268 216 269 217
rect 269 216 270 217
rect 270 216 271 217
rect 271 216 272 217
rect 272 216 273 217
rect 273 216 274 217
rect 274 216 275 217
rect 275 216 276 217
rect 276 216 277 217
rect 277 216 278 217
rect 278 216 279 217
rect 279 216 280 217
rect 280 216 281 217
rect 281 216 282 217
rect 282 216 283 217
rect 283 216 284 217
rect 284 216 285 217
rect 285 216 286 217
rect 286 216 287 217
rect 287 216 288 217
rect 288 216 289 217
rect 334 216 335 217
rect 335 216 336 217
rect 336 216 337 217
rect 337 216 338 217
rect 338 216 339 217
rect 339 216 340 217
rect 362 216 363 217
rect 363 216 364 217
rect 364 216 365 217
rect 365 216 366 217
rect 366 216 367 217
rect 367 216 368 217
rect 368 216 369 217
rect 106 215 107 216
rect 107 215 108 216
rect 108 215 109 216
rect 109 215 110 216
rect 110 215 111 216
rect 111 215 112 216
rect 112 215 113 216
rect 113 215 114 216
rect 114 215 115 216
rect 115 215 116 216
rect 116 215 117 216
rect 117 215 118 216
rect 118 215 119 216
rect 119 215 120 216
rect 120 215 121 216
rect 121 215 122 216
rect 122 215 123 216
rect 123 215 124 216
rect 124 215 125 216
rect 125 215 126 216
rect 126 215 127 216
rect 127 215 128 216
rect 128 215 129 216
rect 129 215 130 216
rect 130 215 131 216
rect 131 215 132 216
rect 132 215 133 216
rect 133 215 134 216
rect 134 215 135 216
rect 135 215 136 216
rect 136 215 137 216
rect 137 215 138 216
rect 138 215 139 216
rect 139 215 140 216
rect 140 215 141 216
rect 141 215 142 216
rect 142 215 143 216
rect 143 215 144 216
rect 144 215 145 216
rect 145 215 146 216
rect 146 215 147 216
rect 163 215 164 216
rect 164 215 165 216
rect 165 215 166 216
rect 166 215 167 216
rect 183 215 184 216
rect 184 215 185 216
rect 185 215 186 216
rect 186 215 187 216
rect 187 215 188 216
rect 188 215 189 216
rect 189 215 190 216
rect 190 215 191 216
rect 191 215 192 216
rect 192 215 193 216
rect 193 215 194 216
rect 194 215 195 216
rect 195 215 196 216
rect 196 215 197 216
rect 197 215 198 216
rect 198 215 199 216
rect 199 215 200 216
rect 250 215 251 216
rect 251 215 252 216
rect 252 215 253 216
rect 253 215 254 216
rect 254 215 255 216
rect 255 215 256 216
rect 256 215 257 216
rect 257 215 258 216
rect 258 215 259 216
rect 259 215 260 216
rect 260 215 261 216
rect 261 215 262 216
rect 262 215 263 216
rect 263 215 264 216
rect 264 215 265 216
rect 265 215 266 216
rect 266 215 267 216
rect 267 215 268 216
rect 268 215 269 216
rect 269 215 270 216
rect 270 215 271 216
rect 271 215 272 216
rect 272 215 273 216
rect 273 215 274 216
rect 274 215 275 216
rect 275 215 276 216
rect 276 215 277 216
rect 277 215 278 216
rect 278 215 279 216
rect 279 215 280 216
rect 280 215 281 216
rect 281 215 282 216
rect 282 215 283 216
rect 283 215 284 216
rect 284 215 285 216
rect 285 215 286 216
rect 286 215 287 216
rect 287 215 288 216
rect 288 215 289 216
rect 289 215 290 216
rect 334 215 335 216
rect 335 215 336 216
rect 336 215 337 216
rect 337 215 338 216
rect 338 215 339 216
rect 339 215 340 216
rect 362 215 363 216
rect 363 215 364 216
rect 364 215 365 216
rect 365 215 366 216
rect 366 215 367 216
rect 367 215 368 216
rect 368 215 369 216
rect 114 214 115 215
rect 115 214 116 215
rect 116 214 117 215
rect 117 214 118 215
rect 118 214 119 215
rect 119 214 120 215
rect 120 214 121 215
rect 121 214 122 215
rect 122 214 123 215
rect 123 214 124 215
rect 124 214 125 215
rect 125 214 126 215
rect 140 214 141 215
rect 141 214 142 215
rect 142 214 143 215
rect 143 214 144 215
rect 144 214 145 215
rect 145 214 146 215
rect 146 214 147 215
rect 163 214 164 215
rect 164 214 165 215
rect 165 214 166 215
rect 166 214 167 215
rect 182 214 183 215
rect 183 214 184 215
rect 184 214 185 215
rect 185 214 186 215
rect 186 214 187 215
rect 187 214 188 215
rect 188 214 189 215
rect 189 214 190 215
rect 190 214 191 215
rect 191 214 192 215
rect 192 214 193 215
rect 193 214 194 215
rect 194 214 195 215
rect 195 214 196 215
rect 196 214 197 215
rect 197 214 198 215
rect 198 214 199 215
rect 199 214 200 215
rect 200 214 201 215
rect 201 214 202 215
rect 202 214 203 215
rect 251 214 252 215
rect 252 214 253 215
rect 253 214 254 215
rect 254 214 255 215
rect 255 214 256 215
rect 256 214 257 215
rect 257 214 258 215
rect 258 214 259 215
rect 259 214 260 215
rect 260 214 261 215
rect 261 214 262 215
rect 262 214 263 215
rect 263 214 264 215
rect 264 214 265 215
rect 265 214 266 215
rect 266 214 267 215
rect 267 214 268 215
rect 268 214 269 215
rect 269 214 270 215
rect 270 214 271 215
rect 271 214 272 215
rect 272 214 273 215
rect 273 214 274 215
rect 274 214 275 215
rect 275 214 276 215
rect 276 214 277 215
rect 277 214 278 215
rect 278 214 279 215
rect 279 214 280 215
rect 280 214 281 215
rect 281 214 282 215
rect 282 214 283 215
rect 283 214 284 215
rect 284 214 285 215
rect 285 214 286 215
rect 286 214 287 215
rect 287 214 288 215
rect 288 214 289 215
rect 289 214 290 215
rect 290 214 291 215
rect 334 214 335 215
rect 335 214 336 215
rect 336 214 337 215
rect 337 214 338 215
rect 338 214 339 215
rect 339 214 340 215
rect 362 214 363 215
rect 363 214 364 215
rect 364 214 365 215
rect 365 214 366 215
rect 366 214 367 215
rect 367 214 368 215
rect 368 214 369 215
rect 369 214 370 215
rect 140 213 141 214
rect 141 213 142 214
rect 142 213 143 214
rect 143 213 144 214
rect 144 213 145 214
rect 145 213 146 214
rect 146 213 147 214
rect 164 213 165 214
rect 165 213 166 214
rect 166 213 167 214
rect 182 213 183 214
rect 183 213 184 214
rect 184 213 185 214
rect 185 213 186 214
rect 186 213 187 214
rect 187 213 188 214
rect 188 213 189 214
rect 189 213 190 214
rect 190 213 191 214
rect 191 213 192 214
rect 192 213 193 214
rect 193 213 194 214
rect 194 213 195 214
rect 195 213 196 214
rect 196 213 197 214
rect 197 213 198 214
rect 198 213 199 214
rect 199 213 200 214
rect 200 213 201 214
rect 201 213 202 214
rect 202 213 203 214
rect 203 213 204 214
rect 204 213 205 214
rect 252 213 253 214
rect 253 213 254 214
rect 254 213 255 214
rect 255 213 256 214
rect 256 213 257 214
rect 257 213 258 214
rect 258 213 259 214
rect 259 213 260 214
rect 260 213 261 214
rect 261 213 262 214
rect 262 213 263 214
rect 263 213 264 214
rect 264 213 265 214
rect 265 213 266 214
rect 266 213 267 214
rect 267 213 268 214
rect 268 213 269 214
rect 269 213 270 214
rect 270 213 271 214
rect 271 213 272 214
rect 272 213 273 214
rect 273 213 274 214
rect 274 213 275 214
rect 275 213 276 214
rect 276 213 277 214
rect 277 213 278 214
rect 278 213 279 214
rect 279 213 280 214
rect 280 213 281 214
rect 281 213 282 214
rect 282 213 283 214
rect 283 213 284 214
rect 284 213 285 214
rect 285 213 286 214
rect 286 213 287 214
rect 287 213 288 214
rect 288 213 289 214
rect 289 213 290 214
rect 290 213 291 214
rect 291 213 292 214
rect 292 213 293 214
rect 334 213 335 214
rect 335 213 336 214
rect 336 213 337 214
rect 337 213 338 214
rect 338 213 339 214
rect 349 213 350 214
rect 350 213 351 214
rect 363 213 364 214
rect 364 213 365 214
rect 365 213 366 214
rect 366 213 367 214
rect 367 213 368 214
rect 368 213 369 214
rect 369 213 370 214
rect 140 212 141 213
rect 141 212 142 213
rect 142 212 143 213
rect 143 212 144 213
rect 144 212 145 213
rect 145 212 146 213
rect 146 212 147 213
rect 164 212 165 213
rect 165 212 166 213
rect 182 212 183 213
rect 183 212 184 213
rect 184 212 185 213
rect 185 212 186 213
rect 186 212 187 213
rect 187 212 188 213
rect 188 212 189 213
rect 189 212 190 213
rect 190 212 191 213
rect 191 212 192 213
rect 192 212 193 213
rect 193 212 194 213
rect 194 212 195 213
rect 195 212 196 213
rect 196 212 197 213
rect 197 212 198 213
rect 198 212 199 213
rect 199 212 200 213
rect 200 212 201 213
rect 201 212 202 213
rect 202 212 203 213
rect 203 212 204 213
rect 204 212 205 213
rect 205 212 206 213
rect 206 212 207 213
rect 252 212 253 213
rect 253 212 254 213
rect 254 212 255 213
rect 255 212 256 213
rect 256 212 257 213
rect 257 212 258 213
rect 258 212 259 213
rect 259 212 260 213
rect 260 212 261 213
rect 261 212 262 213
rect 262 212 263 213
rect 263 212 264 213
rect 264 212 265 213
rect 265 212 266 213
rect 266 212 267 213
rect 267 212 268 213
rect 268 212 269 213
rect 269 212 270 213
rect 270 212 271 213
rect 271 212 272 213
rect 272 212 273 213
rect 273 212 274 213
rect 274 212 275 213
rect 275 212 276 213
rect 276 212 277 213
rect 277 212 278 213
rect 278 212 279 213
rect 279 212 280 213
rect 280 212 281 213
rect 281 212 282 213
rect 282 212 283 213
rect 283 212 284 213
rect 284 212 285 213
rect 285 212 286 213
rect 286 212 287 213
rect 287 212 288 213
rect 288 212 289 213
rect 289 212 290 213
rect 290 212 291 213
rect 291 212 292 213
rect 292 212 293 213
rect 293 212 294 213
rect 334 212 335 213
rect 335 212 336 213
rect 336 212 337 213
rect 337 212 338 213
rect 338 212 339 213
rect 350 212 351 213
rect 351 212 352 213
rect 352 212 353 213
rect 353 212 354 213
rect 363 212 364 213
rect 364 212 365 213
rect 365 212 366 213
rect 366 212 367 213
rect 367 212 368 213
rect 368 212 369 213
rect 369 212 370 213
rect 140 211 141 212
rect 141 211 142 212
rect 142 211 143 212
rect 143 211 144 212
rect 144 211 145 212
rect 145 211 146 212
rect 146 211 147 212
rect 164 211 165 212
rect 165 211 166 212
rect 182 211 183 212
rect 183 211 184 212
rect 184 211 185 212
rect 185 211 186 212
rect 186 211 187 212
rect 196 211 197 212
rect 197 211 198 212
rect 198 211 199 212
rect 199 211 200 212
rect 200 211 201 212
rect 201 211 202 212
rect 202 211 203 212
rect 203 211 204 212
rect 204 211 205 212
rect 205 211 206 212
rect 206 211 207 212
rect 207 211 208 212
rect 253 211 254 212
rect 254 211 255 212
rect 255 211 256 212
rect 256 211 257 212
rect 257 211 258 212
rect 258 211 259 212
rect 259 211 260 212
rect 260 211 261 212
rect 261 211 262 212
rect 262 211 263 212
rect 263 211 264 212
rect 264 211 265 212
rect 265 211 266 212
rect 266 211 267 212
rect 267 211 268 212
rect 268 211 269 212
rect 269 211 270 212
rect 270 211 271 212
rect 271 211 272 212
rect 272 211 273 212
rect 273 211 274 212
rect 274 211 275 212
rect 275 211 276 212
rect 276 211 277 212
rect 277 211 278 212
rect 278 211 279 212
rect 279 211 280 212
rect 280 211 281 212
rect 281 211 282 212
rect 282 211 283 212
rect 283 211 284 212
rect 284 211 285 212
rect 285 211 286 212
rect 286 211 287 212
rect 287 211 288 212
rect 288 211 289 212
rect 289 211 290 212
rect 290 211 291 212
rect 291 211 292 212
rect 292 211 293 212
rect 293 211 294 212
rect 294 211 295 212
rect 334 211 335 212
rect 335 211 336 212
rect 336 211 337 212
rect 337 211 338 212
rect 338 211 339 212
rect 351 211 352 212
rect 352 211 353 212
rect 353 211 354 212
rect 354 211 355 212
rect 355 211 356 212
rect 363 211 364 212
rect 364 211 365 212
rect 365 211 366 212
rect 366 211 367 212
rect 367 211 368 212
rect 368 211 369 212
rect 369 211 370 212
rect 140 210 141 211
rect 141 210 142 211
rect 142 210 143 211
rect 143 210 144 211
rect 144 210 145 211
rect 145 210 146 211
rect 146 210 147 211
rect 165 210 166 211
rect 183 210 184 211
rect 184 210 185 211
rect 200 210 201 211
rect 201 210 202 211
rect 202 210 203 211
rect 203 210 204 211
rect 204 210 205 211
rect 205 210 206 211
rect 206 210 207 211
rect 207 210 208 211
rect 208 210 209 211
rect 254 210 255 211
rect 255 210 256 211
rect 256 210 257 211
rect 257 210 258 211
rect 258 210 259 211
rect 259 210 260 211
rect 260 210 261 211
rect 261 210 262 211
rect 262 210 263 211
rect 263 210 264 211
rect 264 210 265 211
rect 265 210 266 211
rect 266 210 267 211
rect 267 210 268 211
rect 268 210 269 211
rect 269 210 270 211
rect 270 210 271 211
rect 271 210 272 211
rect 272 210 273 211
rect 273 210 274 211
rect 274 210 275 211
rect 275 210 276 211
rect 276 210 277 211
rect 277 210 278 211
rect 278 210 279 211
rect 279 210 280 211
rect 280 210 281 211
rect 281 210 282 211
rect 282 210 283 211
rect 283 210 284 211
rect 284 210 285 211
rect 285 210 286 211
rect 286 210 287 211
rect 287 210 288 211
rect 288 210 289 211
rect 289 210 290 211
rect 290 210 291 211
rect 291 210 292 211
rect 292 210 293 211
rect 293 210 294 211
rect 294 210 295 211
rect 295 210 296 211
rect 333 210 334 211
rect 334 210 335 211
rect 335 210 336 211
rect 336 210 337 211
rect 337 210 338 211
rect 338 210 339 211
rect 352 210 353 211
rect 353 210 354 211
rect 354 210 355 211
rect 355 210 356 211
rect 356 210 357 211
rect 357 210 358 211
rect 363 210 364 211
rect 364 210 365 211
rect 365 210 366 211
rect 366 210 367 211
rect 367 210 368 211
rect 368 210 369 211
rect 369 210 370 211
rect 140 209 141 210
rect 141 209 142 210
rect 142 209 143 210
rect 143 209 144 210
rect 144 209 145 210
rect 145 209 146 210
rect 146 209 147 210
rect 183 209 184 210
rect 203 209 204 210
rect 204 209 205 210
rect 205 209 206 210
rect 206 209 207 210
rect 207 209 208 210
rect 208 209 209 210
rect 209 209 210 210
rect 255 209 256 210
rect 256 209 257 210
rect 257 209 258 210
rect 258 209 259 210
rect 259 209 260 210
rect 260 209 261 210
rect 261 209 262 210
rect 262 209 263 210
rect 263 209 264 210
rect 264 209 265 210
rect 265 209 266 210
rect 266 209 267 210
rect 267 209 268 210
rect 268 209 269 210
rect 269 209 270 210
rect 270 209 271 210
rect 271 209 272 210
rect 272 209 273 210
rect 273 209 274 210
rect 274 209 275 210
rect 275 209 276 210
rect 276 209 277 210
rect 277 209 278 210
rect 278 209 279 210
rect 279 209 280 210
rect 280 209 281 210
rect 281 209 282 210
rect 282 209 283 210
rect 283 209 284 210
rect 284 209 285 210
rect 285 209 286 210
rect 286 209 287 210
rect 287 209 288 210
rect 288 209 289 210
rect 289 209 290 210
rect 290 209 291 210
rect 291 209 292 210
rect 292 209 293 210
rect 293 209 294 210
rect 294 209 295 210
rect 295 209 296 210
rect 296 209 297 210
rect 297 209 298 210
rect 333 209 334 210
rect 334 209 335 210
rect 335 209 336 210
rect 336 209 337 210
rect 337 209 338 210
rect 338 209 339 210
rect 353 209 354 210
rect 354 209 355 210
rect 355 209 356 210
rect 356 209 357 210
rect 357 209 358 210
rect 358 209 359 210
rect 363 209 364 210
rect 364 209 365 210
rect 365 209 366 210
rect 366 209 367 210
rect 367 209 368 210
rect 368 209 369 210
rect 369 209 370 210
rect 140 208 141 209
rect 141 208 142 209
rect 142 208 143 209
rect 143 208 144 209
rect 144 208 145 209
rect 145 208 146 209
rect 146 208 147 209
rect 205 208 206 209
rect 206 208 207 209
rect 207 208 208 209
rect 208 208 209 209
rect 209 208 210 209
rect 210 208 211 209
rect 256 208 257 209
rect 257 208 258 209
rect 258 208 259 209
rect 259 208 260 209
rect 260 208 261 209
rect 261 208 262 209
rect 262 208 263 209
rect 263 208 264 209
rect 264 208 265 209
rect 265 208 266 209
rect 266 208 267 209
rect 267 208 268 209
rect 268 208 269 209
rect 269 208 270 209
rect 270 208 271 209
rect 271 208 272 209
rect 272 208 273 209
rect 273 208 274 209
rect 274 208 275 209
rect 275 208 276 209
rect 276 208 277 209
rect 277 208 278 209
rect 278 208 279 209
rect 279 208 280 209
rect 280 208 281 209
rect 281 208 282 209
rect 282 208 283 209
rect 283 208 284 209
rect 284 208 285 209
rect 285 208 286 209
rect 286 208 287 209
rect 287 208 288 209
rect 288 208 289 209
rect 289 208 290 209
rect 290 208 291 209
rect 291 208 292 209
rect 292 208 293 209
rect 293 208 294 209
rect 294 208 295 209
rect 295 208 296 209
rect 296 208 297 209
rect 297 208 298 209
rect 298 208 299 209
rect 333 208 334 209
rect 334 208 335 209
rect 335 208 336 209
rect 336 208 337 209
rect 337 208 338 209
rect 338 208 339 209
rect 354 208 355 209
rect 355 208 356 209
rect 356 208 357 209
rect 357 208 358 209
rect 358 208 359 209
rect 359 208 360 209
rect 364 208 365 209
rect 365 208 366 209
rect 366 208 367 209
rect 367 208 368 209
rect 368 208 369 209
rect 369 208 370 209
rect 140 207 141 208
rect 141 207 142 208
rect 142 207 143 208
rect 143 207 144 208
rect 144 207 145 208
rect 145 207 146 208
rect 146 207 147 208
rect 207 207 208 208
rect 208 207 209 208
rect 209 207 210 208
rect 210 207 211 208
rect 211 207 212 208
rect 256 207 257 208
rect 257 207 258 208
rect 258 207 259 208
rect 259 207 260 208
rect 260 207 261 208
rect 261 207 262 208
rect 262 207 263 208
rect 263 207 264 208
rect 264 207 265 208
rect 265 207 266 208
rect 266 207 267 208
rect 267 207 268 208
rect 268 207 269 208
rect 269 207 270 208
rect 270 207 271 208
rect 271 207 272 208
rect 272 207 273 208
rect 273 207 274 208
rect 274 207 275 208
rect 275 207 276 208
rect 276 207 277 208
rect 277 207 278 208
rect 278 207 279 208
rect 279 207 280 208
rect 280 207 281 208
rect 281 207 282 208
rect 282 207 283 208
rect 283 207 284 208
rect 284 207 285 208
rect 285 207 286 208
rect 286 207 287 208
rect 287 207 288 208
rect 288 207 289 208
rect 289 207 290 208
rect 290 207 291 208
rect 291 207 292 208
rect 292 207 293 208
rect 293 207 294 208
rect 294 207 295 208
rect 295 207 296 208
rect 296 207 297 208
rect 297 207 298 208
rect 298 207 299 208
rect 299 207 300 208
rect 300 207 301 208
rect 333 207 334 208
rect 334 207 335 208
rect 335 207 336 208
rect 336 207 337 208
rect 337 207 338 208
rect 338 207 339 208
rect 355 207 356 208
rect 356 207 357 208
rect 357 207 358 208
rect 358 207 359 208
rect 359 207 360 208
rect 360 207 361 208
rect 364 207 365 208
rect 365 207 366 208
rect 366 207 367 208
rect 367 207 368 208
rect 368 207 369 208
rect 369 207 370 208
rect 139 206 140 207
rect 140 206 141 207
rect 141 206 142 207
rect 142 206 143 207
rect 143 206 144 207
rect 144 206 145 207
rect 145 206 146 207
rect 146 206 147 207
rect 208 206 209 207
rect 209 206 210 207
rect 210 206 211 207
rect 211 206 212 207
rect 257 206 258 207
rect 258 206 259 207
rect 259 206 260 207
rect 260 206 261 207
rect 261 206 262 207
rect 262 206 263 207
rect 263 206 264 207
rect 264 206 265 207
rect 265 206 266 207
rect 266 206 267 207
rect 267 206 268 207
rect 268 206 269 207
rect 269 206 270 207
rect 270 206 271 207
rect 271 206 272 207
rect 272 206 273 207
rect 273 206 274 207
rect 274 206 275 207
rect 275 206 276 207
rect 276 206 277 207
rect 277 206 278 207
rect 278 206 279 207
rect 279 206 280 207
rect 280 206 281 207
rect 281 206 282 207
rect 282 206 283 207
rect 283 206 284 207
rect 284 206 285 207
rect 285 206 286 207
rect 286 206 287 207
rect 287 206 288 207
rect 290 206 291 207
rect 291 206 292 207
rect 292 206 293 207
rect 293 206 294 207
rect 294 206 295 207
rect 295 206 296 207
rect 296 206 297 207
rect 297 206 298 207
rect 298 206 299 207
rect 299 206 300 207
rect 300 206 301 207
rect 301 206 302 207
rect 302 206 303 207
rect 332 206 333 207
rect 333 206 334 207
rect 334 206 335 207
rect 335 206 336 207
rect 336 206 337 207
rect 337 206 338 207
rect 338 206 339 207
rect 356 206 357 207
rect 357 206 358 207
rect 358 206 359 207
rect 359 206 360 207
rect 360 206 361 207
rect 361 206 362 207
rect 363 206 364 207
rect 364 206 365 207
rect 365 206 366 207
rect 366 206 367 207
rect 367 206 368 207
rect 368 206 369 207
rect 369 206 370 207
rect 139 205 140 206
rect 140 205 141 206
rect 141 205 142 206
rect 142 205 143 206
rect 143 205 144 206
rect 144 205 145 206
rect 145 205 146 206
rect 210 205 211 206
rect 211 205 212 206
rect 258 205 259 206
rect 259 205 260 206
rect 260 205 261 206
rect 261 205 262 206
rect 262 205 263 206
rect 263 205 264 206
rect 264 205 265 206
rect 265 205 266 206
rect 266 205 267 206
rect 267 205 268 206
rect 268 205 269 206
rect 269 205 270 206
rect 270 205 271 206
rect 271 205 272 206
rect 272 205 273 206
rect 273 205 274 206
rect 274 205 275 206
rect 275 205 276 206
rect 276 205 277 206
rect 277 205 278 206
rect 278 205 279 206
rect 279 205 280 206
rect 280 205 281 206
rect 281 205 282 206
rect 282 205 283 206
rect 283 205 284 206
rect 284 205 285 206
rect 285 205 286 206
rect 286 205 287 206
rect 287 205 288 206
rect 292 205 293 206
rect 293 205 294 206
rect 294 205 295 206
rect 295 205 296 206
rect 296 205 297 206
rect 297 205 298 206
rect 298 205 299 206
rect 299 205 300 206
rect 300 205 301 206
rect 301 205 302 206
rect 302 205 303 206
rect 303 205 304 206
rect 304 205 305 206
rect 332 205 333 206
rect 333 205 334 206
rect 334 205 335 206
rect 335 205 336 206
rect 336 205 337 206
rect 337 205 338 206
rect 338 205 339 206
rect 356 205 357 206
rect 357 205 358 206
rect 358 205 359 206
rect 359 205 360 206
rect 360 205 361 206
rect 361 205 362 206
rect 363 205 364 206
rect 364 205 365 206
rect 365 205 366 206
rect 366 205 367 206
rect 367 205 368 206
rect 368 205 369 206
rect 369 205 370 206
rect 139 204 140 205
rect 140 204 141 205
rect 141 204 142 205
rect 142 204 143 205
rect 143 204 144 205
rect 144 204 145 205
rect 145 204 146 205
rect 211 204 212 205
rect 212 204 213 205
rect 259 204 260 205
rect 260 204 261 205
rect 261 204 262 205
rect 262 204 263 205
rect 263 204 264 205
rect 264 204 265 205
rect 265 204 266 205
rect 266 204 267 205
rect 267 204 268 205
rect 268 204 269 205
rect 269 204 270 205
rect 270 204 271 205
rect 271 204 272 205
rect 272 204 273 205
rect 273 204 274 205
rect 274 204 275 205
rect 275 204 276 205
rect 276 204 277 205
rect 277 204 278 205
rect 278 204 279 205
rect 279 204 280 205
rect 280 204 281 205
rect 281 204 282 205
rect 282 204 283 205
rect 283 204 284 205
rect 284 204 285 205
rect 285 204 286 205
rect 286 204 287 205
rect 287 204 288 205
rect 288 204 289 205
rect 289 204 290 205
rect 294 204 295 205
rect 295 204 296 205
rect 296 204 297 205
rect 297 204 298 205
rect 298 204 299 205
rect 299 204 300 205
rect 300 204 301 205
rect 301 204 302 205
rect 302 204 303 205
rect 303 204 304 205
rect 304 204 305 205
rect 305 204 306 205
rect 332 204 333 205
rect 333 204 334 205
rect 334 204 335 205
rect 335 204 336 205
rect 336 204 337 205
rect 337 204 338 205
rect 357 204 358 205
rect 358 204 359 205
rect 359 204 360 205
rect 360 204 361 205
rect 361 204 362 205
rect 362 204 363 205
rect 363 204 364 205
rect 364 204 365 205
rect 365 204 366 205
rect 366 204 367 205
rect 367 204 368 205
rect 368 204 369 205
rect 369 204 370 205
rect 139 203 140 204
rect 140 203 141 204
rect 141 203 142 204
rect 142 203 143 204
rect 143 203 144 204
rect 144 203 145 204
rect 145 203 146 204
rect 212 203 213 204
rect 260 203 261 204
rect 261 203 262 204
rect 262 203 263 204
rect 263 203 264 204
rect 264 203 265 204
rect 265 203 266 204
rect 266 203 267 204
rect 267 203 268 204
rect 268 203 269 204
rect 269 203 270 204
rect 270 203 271 204
rect 271 203 272 204
rect 272 203 273 204
rect 273 203 274 204
rect 274 203 275 204
rect 275 203 276 204
rect 276 203 277 204
rect 277 203 278 204
rect 278 203 279 204
rect 279 203 280 204
rect 280 203 281 204
rect 281 203 282 204
rect 282 203 283 204
rect 283 203 284 204
rect 284 203 285 204
rect 285 203 286 204
rect 286 203 287 204
rect 287 203 288 204
rect 288 203 289 204
rect 289 203 290 204
rect 290 203 291 204
rect 297 203 298 204
rect 298 203 299 204
rect 299 203 300 204
rect 300 203 301 204
rect 301 203 302 204
rect 302 203 303 204
rect 331 203 332 204
rect 332 203 333 204
rect 333 203 334 204
rect 334 203 335 204
rect 335 203 336 204
rect 336 203 337 204
rect 337 203 338 204
rect 357 203 358 204
rect 358 203 359 204
rect 359 203 360 204
rect 360 203 361 204
rect 361 203 362 204
rect 362 203 363 204
rect 363 203 364 204
rect 364 203 365 204
rect 365 203 366 204
rect 366 203 367 204
rect 367 203 368 204
rect 368 203 369 204
rect 138 202 139 203
rect 139 202 140 203
rect 140 202 141 203
rect 141 202 142 203
rect 142 202 143 203
rect 143 202 144 203
rect 144 202 145 203
rect 260 202 261 203
rect 261 202 262 203
rect 262 202 263 203
rect 263 202 264 203
rect 264 202 265 203
rect 265 202 266 203
rect 266 202 267 203
rect 267 202 268 203
rect 269 202 270 203
rect 270 202 271 203
rect 271 202 272 203
rect 272 202 273 203
rect 273 202 274 203
rect 274 202 275 203
rect 275 202 276 203
rect 276 202 277 203
rect 277 202 278 203
rect 278 202 279 203
rect 279 202 280 203
rect 280 202 281 203
rect 281 202 282 203
rect 282 202 283 203
rect 283 202 284 203
rect 284 202 285 203
rect 285 202 286 203
rect 286 202 287 203
rect 287 202 288 203
rect 288 202 289 203
rect 289 202 290 203
rect 290 202 291 203
rect 291 202 292 203
rect 292 202 293 203
rect 331 202 332 203
rect 332 202 333 203
rect 333 202 334 203
rect 334 202 335 203
rect 335 202 336 203
rect 336 202 337 203
rect 337 202 338 203
rect 358 202 359 203
rect 359 202 360 203
rect 360 202 361 203
rect 361 202 362 203
rect 362 202 363 203
rect 363 202 364 203
rect 364 202 365 203
rect 365 202 366 203
rect 366 202 367 203
rect 367 202 368 203
rect 368 202 369 203
rect 138 201 139 202
rect 139 201 140 202
rect 140 201 141 202
rect 141 201 142 202
rect 142 201 143 202
rect 143 201 144 202
rect 144 201 145 202
rect 261 201 262 202
rect 262 201 263 202
rect 263 201 264 202
rect 264 201 265 202
rect 265 201 266 202
rect 266 201 267 202
rect 267 201 268 202
rect 271 201 272 202
rect 272 201 273 202
rect 273 201 274 202
rect 274 201 275 202
rect 275 201 276 202
rect 276 201 277 202
rect 277 201 278 202
rect 278 201 279 202
rect 279 201 280 202
rect 280 201 281 202
rect 281 201 282 202
rect 282 201 283 202
rect 283 201 284 202
rect 284 201 285 202
rect 285 201 286 202
rect 286 201 287 202
rect 287 201 288 202
rect 288 201 289 202
rect 289 201 290 202
rect 290 201 291 202
rect 291 201 292 202
rect 292 201 293 202
rect 293 201 294 202
rect 294 201 295 202
rect 295 201 296 202
rect 330 201 331 202
rect 331 201 332 202
rect 332 201 333 202
rect 333 201 334 202
rect 334 201 335 202
rect 335 201 336 202
rect 336 201 337 202
rect 337 201 338 202
rect 358 201 359 202
rect 359 201 360 202
rect 360 201 361 202
rect 361 201 362 202
rect 362 201 363 202
rect 363 201 364 202
rect 364 201 365 202
rect 365 201 366 202
rect 366 201 367 202
rect 367 201 368 202
rect 368 201 369 202
rect 137 200 138 201
rect 138 200 139 201
rect 139 200 140 201
rect 140 200 141 201
rect 141 200 142 201
rect 142 200 143 201
rect 143 200 144 201
rect 144 200 145 201
rect 262 200 263 201
rect 263 200 264 201
rect 264 200 265 201
rect 265 200 266 201
rect 266 200 267 201
rect 267 200 268 201
rect 274 200 275 201
rect 275 200 276 201
rect 276 200 277 201
rect 277 200 278 201
rect 278 200 279 201
rect 279 200 280 201
rect 280 200 281 201
rect 281 200 282 201
rect 282 200 283 201
rect 283 200 284 201
rect 284 200 285 201
rect 285 200 286 201
rect 286 200 287 201
rect 287 200 288 201
rect 288 200 289 201
rect 289 200 290 201
rect 290 200 291 201
rect 291 200 292 201
rect 292 200 293 201
rect 293 200 294 201
rect 294 200 295 201
rect 295 200 296 201
rect 296 200 297 201
rect 297 200 298 201
rect 330 200 331 201
rect 331 200 332 201
rect 332 200 333 201
rect 333 200 334 201
rect 334 200 335 201
rect 335 200 336 201
rect 336 200 337 201
rect 337 200 338 201
rect 358 200 359 201
rect 359 200 360 201
rect 360 200 361 201
rect 361 200 362 201
rect 362 200 363 201
rect 363 200 364 201
rect 364 200 365 201
rect 365 200 366 201
rect 366 200 367 201
rect 367 200 368 201
rect 136 199 137 200
rect 137 199 138 200
rect 138 199 139 200
rect 139 199 140 200
rect 140 199 141 200
rect 141 199 142 200
rect 142 199 143 200
rect 143 199 144 200
rect 263 199 264 200
rect 264 199 265 200
rect 265 199 266 200
rect 266 199 267 200
rect 267 199 268 200
rect 268 199 269 200
rect 276 199 277 200
rect 277 199 278 200
rect 278 199 279 200
rect 279 199 280 200
rect 280 199 281 200
rect 281 199 282 200
rect 282 199 283 200
rect 283 199 284 200
rect 284 199 285 200
rect 285 199 286 200
rect 286 199 287 200
rect 287 199 288 200
rect 288 199 289 200
rect 289 199 290 200
rect 290 199 291 200
rect 291 199 292 200
rect 292 199 293 200
rect 293 199 294 200
rect 294 199 295 200
rect 295 199 296 200
rect 296 199 297 200
rect 297 199 298 200
rect 298 199 299 200
rect 299 199 300 200
rect 329 199 330 200
rect 330 199 331 200
rect 331 199 332 200
rect 332 199 333 200
rect 333 199 334 200
rect 334 199 335 200
rect 335 199 336 200
rect 336 199 337 200
rect 359 199 360 200
rect 360 199 361 200
rect 361 199 362 200
rect 362 199 363 200
rect 363 199 364 200
rect 364 199 365 200
rect 365 199 366 200
rect 366 199 367 200
rect 367 199 368 200
rect 136 198 137 199
rect 137 198 138 199
rect 138 198 139 199
rect 139 198 140 199
rect 140 198 141 199
rect 141 198 142 199
rect 142 198 143 199
rect 143 198 144 199
rect 263 198 264 199
rect 264 198 265 199
rect 265 198 266 199
rect 266 198 267 199
rect 267 198 268 199
rect 268 198 269 199
rect 280 198 281 199
rect 281 198 282 199
rect 282 198 283 199
rect 283 198 284 199
rect 284 198 285 199
rect 285 198 286 199
rect 286 198 287 199
rect 287 198 288 199
rect 288 198 289 199
rect 289 198 290 199
rect 290 198 291 199
rect 291 198 292 199
rect 292 198 293 199
rect 293 198 294 199
rect 294 198 295 199
rect 295 198 296 199
rect 296 198 297 199
rect 329 198 330 199
rect 330 198 331 199
rect 331 198 332 199
rect 332 198 333 199
rect 333 198 334 199
rect 334 198 335 199
rect 335 198 336 199
rect 336 198 337 199
rect 337 198 338 199
rect 338 198 339 199
rect 339 198 340 199
rect 359 198 360 199
rect 360 198 361 199
rect 361 198 362 199
rect 362 198 363 199
rect 363 198 364 199
rect 364 198 365 199
rect 365 198 366 199
rect 366 198 367 199
rect 135 197 136 198
rect 136 197 137 198
rect 137 197 138 198
rect 138 197 139 198
rect 139 197 140 198
rect 140 197 141 198
rect 141 197 142 198
rect 142 197 143 198
rect 264 197 265 198
rect 265 197 266 198
rect 266 197 267 198
rect 267 197 268 198
rect 268 197 269 198
rect 287 197 288 198
rect 288 197 289 198
rect 289 197 290 198
rect 290 197 291 198
rect 328 197 329 198
rect 329 197 330 198
rect 330 197 331 198
rect 331 197 332 198
rect 332 197 333 198
rect 333 197 334 198
rect 334 197 335 198
rect 335 197 336 198
rect 336 197 337 198
rect 337 197 338 198
rect 338 197 339 198
rect 339 197 340 198
rect 340 197 341 198
rect 341 197 342 198
rect 359 197 360 198
rect 360 197 361 198
rect 361 197 362 198
rect 362 197 363 198
rect 363 197 364 198
rect 364 197 365 198
rect 365 197 366 198
rect 135 196 136 197
rect 136 196 137 197
rect 137 196 138 197
rect 138 196 139 197
rect 139 196 140 197
rect 140 196 141 197
rect 141 196 142 197
rect 142 196 143 197
rect 265 196 266 197
rect 266 196 267 197
rect 267 196 268 197
rect 268 196 269 197
rect 269 196 270 197
rect 327 196 328 197
rect 328 196 329 197
rect 329 196 330 197
rect 330 196 331 197
rect 331 196 332 197
rect 332 196 333 197
rect 333 196 334 197
rect 334 196 335 197
rect 335 196 336 197
rect 336 196 337 197
rect 337 196 338 197
rect 338 196 339 197
rect 339 196 340 197
rect 340 196 341 197
rect 341 196 342 197
rect 342 196 343 197
rect 343 196 344 197
rect 359 196 360 197
rect 360 196 361 197
rect 361 196 362 197
rect 362 196 363 197
rect 363 196 364 197
rect 364 196 365 197
rect 365 196 366 197
rect 134 195 135 196
rect 135 195 136 196
rect 136 195 137 196
rect 137 195 138 196
rect 138 195 139 196
rect 139 195 140 196
rect 140 195 141 196
rect 141 195 142 196
rect 142 195 143 196
rect 265 195 266 196
rect 266 195 267 196
rect 267 195 268 196
rect 268 195 269 196
rect 269 195 270 196
rect 327 195 328 196
rect 328 195 329 196
rect 329 195 330 196
rect 330 195 331 196
rect 331 195 332 196
rect 332 195 333 196
rect 333 195 334 196
rect 334 195 335 196
rect 335 195 336 196
rect 336 195 337 196
rect 337 195 338 196
rect 338 195 339 196
rect 339 195 340 196
rect 340 195 341 196
rect 341 195 342 196
rect 342 195 343 196
rect 343 195 344 196
rect 344 195 345 196
rect 359 195 360 196
rect 360 195 361 196
rect 361 195 362 196
rect 362 195 363 196
rect 363 195 364 196
rect 364 195 365 196
rect 365 195 366 196
rect 134 194 135 195
rect 135 194 136 195
rect 136 194 137 195
rect 137 194 138 195
rect 138 194 139 195
rect 139 194 140 195
rect 140 194 141 195
rect 141 194 142 195
rect 266 194 267 195
rect 267 194 268 195
rect 268 194 269 195
rect 269 194 270 195
rect 270 194 271 195
rect 326 194 327 195
rect 327 194 328 195
rect 328 194 329 195
rect 329 194 330 195
rect 330 194 331 195
rect 331 194 332 195
rect 332 194 333 195
rect 333 194 334 195
rect 334 194 335 195
rect 337 194 338 195
rect 338 194 339 195
rect 339 194 340 195
rect 340 194 341 195
rect 341 194 342 195
rect 342 194 343 195
rect 343 194 344 195
rect 344 194 345 195
rect 345 194 346 195
rect 359 194 360 195
rect 360 194 361 195
rect 361 194 362 195
rect 362 194 363 195
rect 363 194 364 195
rect 364 194 365 195
rect 365 194 366 195
rect 133 193 134 194
rect 134 193 135 194
rect 135 193 136 194
rect 136 193 137 194
rect 137 193 138 194
rect 138 193 139 194
rect 139 193 140 194
rect 140 193 141 194
rect 141 193 142 194
rect 267 193 268 194
rect 268 193 269 194
rect 269 193 270 194
rect 270 193 271 194
rect 325 193 326 194
rect 326 193 327 194
rect 327 193 328 194
rect 328 193 329 194
rect 329 193 330 194
rect 330 193 331 194
rect 331 193 332 194
rect 332 193 333 194
rect 333 193 334 194
rect 334 193 335 194
rect 337 193 338 194
rect 338 193 339 194
rect 339 193 340 194
rect 340 193 341 194
rect 341 193 342 194
rect 342 193 343 194
rect 343 193 344 194
rect 344 193 345 194
rect 345 193 346 194
rect 346 193 347 194
rect 359 193 360 194
rect 360 193 361 194
rect 361 193 362 194
rect 362 193 363 194
rect 363 193 364 194
rect 364 193 365 194
rect 365 193 366 194
rect 133 192 134 193
rect 134 192 135 193
rect 135 192 136 193
rect 136 192 137 193
rect 137 192 138 193
rect 138 192 139 193
rect 139 192 140 193
rect 140 192 141 193
rect 267 192 268 193
rect 268 192 269 193
rect 269 192 270 193
rect 270 192 271 193
rect 271 192 272 193
rect 325 192 326 193
rect 326 192 327 193
rect 327 192 328 193
rect 328 192 329 193
rect 329 192 330 193
rect 330 192 331 193
rect 331 192 332 193
rect 332 192 333 193
rect 333 192 334 193
rect 337 192 338 193
rect 338 192 339 193
rect 339 192 340 193
rect 340 192 341 193
rect 341 192 342 193
rect 342 192 343 193
rect 343 192 344 193
rect 344 192 345 193
rect 345 192 346 193
rect 346 192 347 193
rect 347 192 348 193
rect 359 192 360 193
rect 360 192 361 193
rect 361 192 362 193
rect 362 192 363 193
rect 363 192 364 193
rect 364 192 365 193
rect 365 192 366 193
rect 132 191 133 192
rect 133 191 134 192
rect 134 191 135 192
rect 135 191 136 192
rect 136 191 137 192
rect 137 191 138 192
rect 138 191 139 192
rect 139 191 140 192
rect 268 191 269 192
rect 269 191 270 192
rect 270 191 271 192
rect 271 191 272 192
rect 324 191 325 192
rect 325 191 326 192
rect 326 191 327 192
rect 327 191 328 192
rect 328 191 329 192
rect 329 191 330 192
rect 330 191 331 192
rect 331 191 332 192
rect 332 191 333 192
rect 337 191 338 192
rect 338 191 339 192
rect 339 191 340 192
rect 340 191 341 192
rect 341 191 342 192
rect 342 191 343 192
rect 343 191 344 192
rect 344 191 345 192
rect 345 191 346 192
rect 346 191 347 192
rect 347 191 348 192
rect 348 191 349 192
rect 358 191 359 192
rect 359 191 360 192
rect 360 191 361 192
rect 361 191 362 192
rect 362 191 363 192
rect 363 191 364 192
rect 364 191 365 192
rect 365 191 366 192
rect 132 190 133 191
rect 133 190 134 191
rect 134 190 135 191
rect 135 190 136 191
rect 136 190 137 191
rect 137 190 138 191
rect 138 190 139 191
rect 139 190 140 191
rect 269 190 270 191
rect 270 190 271 191
rect 271 190 272 191
rect 323 190 324 191
rect 324 190 325 191
rect 325 190 326 191
rect 326 190 327 191
rect 327 190 328 191
rect 328 190 329 191
rect 329 190 330 191
rect 330 190 331 191
rect 331 190 332 191
rect 332 190 333 191
rect 337 190 338 191
rect 338 190 339 191
rect 339 190 340 191
rect 340 190 341 191
rect 341 190 342 191
rect 342 190 343 191
rect 343 190 344 191
rect 344 190 345 191
rect 345 190 346 191
rect 346 190 347 191
rect 347 190 348 191
rect 348 190 349 191
rect 349 190 350 191
rect 358 190 359 191
rect 359 190 360 191
rect 360 190 361 191
rect 361 190 362 191
rect 362 190 363 191
rect 363 190 364 191
rect 364 190 365 191
rect 131 189 132 190
rect 132 189 133 190
rect 133 189 134 190
rect 134 189 135 190
rect 135 189 136 190
rect 136 189 137 190
rect 137 189 138 190
rect 138 189 139 190
rect 139 189 140 190
rect 270 189 271 190
rect 271 189 272 190
rect 272 189 273 190
rect 322 189 323 190
rect 323 189 324 190
rect 324 189 325 190
rect 325 189 326 190
rect 326 189 327 190
rect 327 189 328 190
rect 328 189 329 190
rect 329 189 330 190
rect 330 189 331 190
rect 331 189 332 190
rect 337 189 338 190
rect 338 189 339 190
rect 339 189 340 190
rect 340 189 341 190
rect 341 189 342 190
rect 344 189 345 190
rect 345 189 346 190
rect 346 189 347 190
rect 347 189 348 190
rect 348 189 349 190
rect 349 189 350 190
rect 358 189 359 190
rect 359 189 360 190
rect 360 189 361 190
rect 361 189 362 190
rect 362 189 363 190
rect 363 189 364 190
rect 364 189 365 190
rect 131 188 132 189
rect 132 188 133 189
rect 133 188 134 189
rect 134 188 135 189
rect 135 188 136 189
rect 136 188 137 189
rect 137 188 138 189
rect 138 188 139 189
rect 139 188 140 189
rect 270 188 271 189
rect 271 188 272 189
rect 272 188 273 189
rect 321 188 322 189
rect 322 188 323 189
rect 323 188 324 189
rect 324 188 325 189
rect 325 188 326 189
rect 326 188 327 189
rect 327 188 328 189
rect 328 188 329 189
rect 329 188 330 189
rect 330 188 331 189
rect 337 188 338 189
rect 338 188 339 189
rect 339 188 340 189
rect 340 188 341 189
rect 345 188 346 189
rect 346 188 347 189
rect 347 188 348 189
rect 348 188 349 189
rect 349 188 350 189
rect 350 188 351 189
rect 358 188 359 189
rect 359 188 360 189
rect 360 188 361 189
rect 361 188 362 189
rect 362 188 363 189
rect 363 188 364 189
rect 364 188 365 189
rect 130 187 131 188
rect 131 187 132 188
rect 132 187 133 188
rect 133 187 134 188
rect 134 187 135 188
rect 135 187 136 188
rect 136 187 137 188
rect 137 187 138 188
rect 138 187 139 188
rect 271 187 272 188
rect 272 187 273 188
rect 320 187 321 188
rect 321 187 322 188
rect 322 187 323 188
rect 323 187 324 188
rect 324 187 325 188
rect 325 187 326 188
rect 326 187 327 188
rect 327 187 328 188
rect 328 187 329 188
rect 329 187 330 188
rect 337 187 338 188
rect 338 187 339 188
rect 339 187 340 188
rect 340 187 341 188
rect 345 187 346 188
rect 346 187 347 188
rect 347 187 348 188
rect 348 187 349 188
rect 349 187 350 188
rect 350 187 351 188
rect 357 187 358 188
rect 358 187 359 188
rect 359 187 360 188
rect 360 187 361 188
rect 361 187 362 188
rect 362 187 363 188
rect 363 187 364 188
rect 364 187 365 188
rect 130 186 131 187
rect 131 186 132 187
rect 132 186 133 187
rect 133 186 134 187
rect 134 186 135 187
rect 135 186 136 187
rect 136 186 137 187
rect 137 186 138 187
rect 138 186 139 187
rect 272 186 273 187
rect 319 186 320 187
rect 320 186 321 187
rect 321 186 322 187
rect 322 186 323 187
rect 323 186 324 187
rect 324 186 325 187
rect 325 186 326 187
rect 326 186 327 187
rect 327 186 328 187
rect 328 186 329 187
rect 329 186 330 187
rect 337 186 338 187
rect 338 186 339 187
rect 339 186 340 187
rect 340 186 341 187
rect 346 186 347 187
rect 347 186 348 187
rect 348 186 349 187
rect 349 186 350 187
rect 350 186 351 187
rect 351 186 352 187
rect 357 186 358 187
rect 358 186 359 187
rect 359 186 360 187
rect 360 186 361 187
rect 361 186 362 187
rect 362 186 363 187
rect 363 186 364 187
rect 130 185 131 186
rect 131 185 132 186
rect 132 185 133 186
rect 133 185 134 186
rect 134 185 135 186
rect 135 185 136 186
rect 136 185 137 186
rect 137 185 138 186
rect 138 185 139 186
rect 272 185 273 186
rect 318 185 319 186
rect 319 185 320 186
rect 320 185 321 186
rect 321 185 322 186
rect 322 185 323 186
rect 323 185 324 186
rect 324 185 325 186
rect 325 185 326 186
rect 326 185 327 186
rect 327 185 328 186
rect 328 185 329 186
rect 337 185 338 186
rect 338 185 339 186
rect 339 185 340 186
rect 340 185 341 186
rect 346 185 347 186
rect 347 185 348 186
rect 348 185 349 186
rect 349 185 350 186
rect 350 185 351 186
rect 351 185 352 186
rect 356 185 357 186
rect 357 185 358 186
rect 358 185 359 186
rect 359 185 360 186
rect 360 185 361 186
rect 361 185 362 186
rect 362 185 363 186
rect 363 185 364 186
rect 130 184 131 185
rect 131 184 132 185
rect 132 184 133 185
rect 133 184 134 185
rect 134 184 135 185
rect 135 184 136 185
rect 136 184 137 185
rect 137 184 138 185
rect 138 184 139 185
rect 317 184 318 185
rect 318 184 319 185
rect 319 184 320 185
rect 320 184 321 185
rect 321 184 322 185
rect 322 184 323 185
rect 323 184 324 185
rect 324 184 325 185
rect 325 184 326 185
rect 326 184 327 185
rect 327 184 328 185
rect 338 184 339 185
rect 339 184 340 185
rect 340 184 341 185
rect 346 184 347 185
rect 347 184 348 185
rect 348 184 349 185
rect 349 184 350 185
rect 350 184 351 185
rect 351 184 352 185
rect 352 184 353 185
rect 356 184 357 185
rect 357 184 358 185
rect 358 184 359 185
rect 359 184 360 185
rect 360 184 361 185
rect 361 184 362 185
rect 362 184 363 185
rect 363 184 364 185
rect 130 183 131 184
rect 131 183 132 184
rect 132 183 133 184
rect 133 183 134 184
rect 134 183 135 184
rect 135 183 136 184
rect 136 183 137 184
rect 137 183 138 184
rect 138 183 139 184
rect 139 183 140 184
rect 315 183 316 184
rect 316 183 317 184
rect 317 183 318 184
rect 318 183 319 184
rect 319 183 320 184
rect 320 183 321 184
rect 321 183 322 184
rect 322 183 323 184
rect 323 183 324 184
rect 324 183 325 184
rect 325 183 326 184
rect 326 183 327 184
rect 338 183 339 184
rect 339 183 340 184
rect 340 183 341 184
rect 347 183 348 184
rect 348 183 349 184
rect 349 183 350 184
rect 350 183 351 184
rect 351 183 352 184
rect 352 183 353 184
rect 355 183 356 184
rect 356 183 357 184
rect 357 183 358 184
rect 358 183 359 184
rect 359 183 360 184
rect 360 183 361 184
rect 361 183 362 184
rect 362 183 363 184
rect 130 182 131 183
rect 131 182 132 183
rect 132 182 133 183
rect 133 182 134 183
rect 134 182 135 183
rect 135 182 136 183
rect 136 182 137 183
rect 137 182 138 183
rect 138 182 139 183
rect 139 182 140 183
rect 314 182 315 183
rect 315 182 316 183
rect 316 182 317 183
rect 317 182 318 183
rect 318 182 319 183
rect 319 182 320 183
rect 320 182 321 183
rect 321 182 322 183
rect 322 182 323 183
rect 323 182 324 183
rect 324 182 325 183
rect 325 182 326 183
rect 338 182 339 183
rect 339 182 340 183
rect 340 182 341 183
rect 347 182 348 183
rect 348 182 349 183
rect 349 182 350 183
rect 350 182 351 183
rect 351 182 352 183
rect 352 182 353 183
rect 354 182 355 183
rect 355 182 356 183
rect 356 182 357 183
rect 357 182 358 183
rect 358 182 359 183
rect 359 182 360 183
rect 360 182 361 183
rect 361 182 362 183
rect 362 182 363 183
rect 130 181 131 182
rect 131 181 132 182
rect 132 181 133 182
rect 133 181 134 182
rect 134 181 135 182
rect 135 181 136 182
rect 136 181 137 182
rect 137 181 138 182
rect 138 181 139 182
rect 139 181 140 182
rect 312 181 313 182
rect 313 181 314 182
rect 314 181 315 182
rect 315 181 316 182
rect 316 181 317 182
rect 317 181 318 182
rect 318 181 319 182
rect 319 181 320 182
rect 320 181 321 182
rect 321 181 322 182
rect 322 181 323 182
rect 323 181 324 182
rect 324 181 325 182
rect 338 181 339 182
rect 339 181 340 182
rect 340 181 341 182
rect 347 181 348 182
rect 348 181 349 182
rect 349 181 350 182
rect 350 181 351 182
rect 351 181 352 182
rect 352 181 353 182
rect 354 181 355 182
rect 355 181 356 182
rect 356 181 357 182
rect 357 181 358 182
rect 358 181 359 182
rect 359 181 360 182
rect 360 181 361 182
rect 361 181 362 182
rect 131 180 132 181
rect 132 180 133 181
rect 133 180 134 181
rect 134 180 135 181
rect 135 180 136 181
rect 136 180 137 181
rect 137 180 138 181
rect 138 180 139 181
rect 139 180 140 181
rect 140 180 141 181
rect 309 180 310 181
rect 310 180 311 181
rect 311 180 312 181
rect 312 180 313 181
rect 313 180 314 181
rect 314 180 315 181
rect 315 180 316 181
rect 316 180 317 181
rect 317 180 318 181
rect 318 180 319 181
rect 319 180 320 181
rect 320 180 321 181
rect 321 180 322 181
rect 322 180 323 181
rect 323 180 324 181
rect 338 180 339 181
rect 339 180 340 181
rect 340 180 341 181
rect 347 180 348 181
rect 348 180 349 181
rect 349 180 350 181
rect 350 180 351 181
rect 351 180 352 181
rect 352 180 353 181
rect 353 180 354 181
rect 354 180 355 181
rect 355 180 356 181
rect 356 180 357 181
rect 357 180 358 181
rect 358 180 359 181
rect 359 180 360 181
rect 360 180 361 181
rect 131 179 132 180
rect 132 179 133 180
rect 133 179 134 180
rect 134 179 135 180
rect 135 179 136 180
rect 136 179 137 180
rect 137 179 138 180
rect 138 179 139 180
rect 139 179 140 180
rect 140 179 141 180
rect 306 179 307 180
rect 307 179 308 180
rect 308 179 309 180
rect 309 179 310 180
rect 310 179 311 180
rect 311 179 312 180
rect 312 179 313 180
rect 313 179 314 180
rect 314 179 315 180
rect 315 179 316 180
rect 316 179 317 180
rect 317 179 318 180
rect 318 179 319 180
rect 319 179 320 180
rect 320 179 321 180
rect 321 179 322 180
rect 322 179 323 180
rect 338 179 339 180
rect 339 179 340 180
rect 348 179 349 180
rect 349 179 350 180
rect 350 179 351 180
rect 351 179 352 180
rect 352 179 353 180
rect 353 179 354 180
rect 354 179 355 180
rect 355 179 356 180
rect 356 179 357 180
rect 357 179 358 180
rect 358 179 359 180
rect 359 179 360 180
rect 360 179 361 180
rect 132 178 133 179
rect 133 178 134 179
rect 134 178 135 179
rect 135 178 136 179
rect 136 178 137 179
rect 137 178 138 179
rect 138 178 139 179
rect 139 178 140 179
rect 140 178 141 179
rect 141 178 142 179
rect 292 178 293 179
rect 293 178 294 179
rect 294 178 295 179
rect 300 178 301 179
rect 301 178 302 179
rect 302 178 303 179
rect 303 178 304 179
rect 304 178 305 179
rect 305 178 306 179
rect 306 178 307 179
rect 307 178 308 179
rect 308 178 309 179
rect 309 178 310 179
rect 310 178 311 179
rect 311 178 312 179
rect 312 178 313 179
rect 313 178 314 179
rect 314 178 315 179
rect 315 178 316 179
rect 316 178 317 179
rect 317 178 318 179
rect 318 178 319 179
rect 319 178 320 179
rect 320 178 321 179
rect 321 178 322 179
rect 338 178 339 179
rect 339 178 340 179
rect 348 178 349 179
rect 349 178 350 179
rect 350 178 351 179
rect 351 178 352 179
rect 352 178 353 179
rect 353 178 354 179
rect 354 178 355 179
rect 355 178 356 179
rect 356 178 357 179
rect 357 178 358 179
rect 358 178 359 179
rect 359 178 360 179
rect 132 177 133 178
rect 133 177 134 178
rect 134 177 135 178
rect 135 177 136 178
rect 136 177 137 178
rect 137 177 138 178
rect 138 177 139 178
rect 139 177 140 178
rect 140 177 141 178
rect 141 177 142 178
rect 291 177 292 178
rect 292 177 293 178
rect 293 177 294 178
rect 294 177 295 178
rect 295 177 296 178
rect 296 177 297 178
rect 297 177 298 178
rect 298 177 299 178
rect 299 177 300 178
rect 300 177 301 178
rect 301 177 302 178
rect 302 177 303 178
rect 303 177 304 178
rect 304 177 305 178
rect 305 177 306 178
rect 306 177 307 178
rect 307 177 308 178
rect 308 177 309 178
rect 309 177 310 178
rect 310 177 311 178
rect 311 177 312 178
rect 312 177 313 178
rect 313 177 314 178
rect 314 177 315 178
rect 315 177 316 178
rect 316 177 317 178
rect 317 177 318 178
rect 318 177 319 178
rect 319 177 320 178
rect 320 177 321 178
rect 338 177 339 178
rect 339 177 340 178
rect 348 177 349 178
rect 349 177 350 178
rect 350 177 351 178
rect 351 177 352 178
rect 352 177 353 178
rect 353 177 354 178
rect 354 177 355 178
rect 355 177 356 178
rect 356 177 357 178
rect 357 177 358 178
rect 358 177 359 178
rect 133 176 134 177
rect 134 176 135 177
rect 135 176 136 177
rect 136 176 137 177
rect 137 176 138 177
rect 138 176 139 177
rect 139 176 140 177
rect 140 176 141 177
rect 141 176 142 177
rect 142 176 143 177
rect 291 176 292 177
rect 292 176 293 177
rect 293 176 294 177
rect 294 176 295 177
rect 295 176 296 177
rect 296 176 297 177
rect 297 176 298 177
rect 298 176 299 177
rect 299 176 300 177
rect 300 176 301 177
rect 301 176 302 177
rect 302 176 303 177
rect 303 176 304 177
rect 304 176 305 177
rect 305 176 306 177
rect 306 176 307 177
rect 307 176 308 177
rect 308 176 309 177
rect 309 176 310 177
rect 310 176 311 177
rect 311 176 312 177
rect 312 176 313 177
rect 313 176 314 177
rect 314 176 315 177
rect 315 176 316 177
rect 316 176 317 177
rect 317 176 318 177
rect 318 176 319 177
rect 338 176 339 177
rect 339 176 340 177
rect 348 176 349 177
rect 349 176 350 177
rect 350 176 351 177
rect 351 176 352 177
rect 352 176 353 177
rect 353 176 354 177
rect 354 176 355 177
rect 355 176 356 177
rect 356 176 357 177
rect 357 176 358 177
rect 133 175 134 176
rect 134 175 135 176
rect 135 175 136 176
rect 136 175 137 176
rect 137 175 138 176
rect 138 175 139 176
rect 139 175 140 176
rect 140 175 141 176
rect 141 175 142 176
rect 142 175 143 176
rect 291 175 292 176
rect 292 175 293 176
rect 293 175 294 176
rect 294 175 295 176
rect 295 175 296 176
rect 296 175 297 176
rect 297 175 298 176
rect 298 175 299 176
rect 299 175 300 176
rect 300 175 301 176
rect 301 175 302 176
rect 302 175 303 176
rect 303 175 304 176
rect 304 175 305 176
rect 305 175 306 176
rect 306 175 307 176
rect 307 175 308 176
rect 308 175 309 176
rect 309 175 310 176
rect 310 175 311 176
rect 311 175 312 176
rect 312 175 313 176
rect 313 175 314 176
rect 314 175 315 176
rect 315 175 316 176
rect 316 175 317 176
rect 317 175 318 176
rect 338 175 339 176
rect 348 175 349 176
rect 349 175 350 176
rect 350 175 351 176
rect 351 175 352 176
rect 352 175 353 176
rect 353 175 354 176
rect 354 175 355 176
rect 355 175 356 176
rect 356 175 357 176
rect 134 174 135 175
rect 135 174 136 175
rect 136 174 137 175
rect 137 174 138 175
rect 138 174 139 175
rect 139 174 140 175
rect 140 174 141 175
rect 141 174 142 175
rect 142 174 143 175
rect 143 174 144 175
rect 290 174 291 175
rect 291 174 292 175
rect 292 174 293 175
rect 293 174 294 175
rect 294 174 295 175
rect 295 174 296 175
rect 296 174 297 175
rect 297 174 298 175
rect 298 174 299 175
rect 299 174 300 175
rect 300 174 301 175
rect 301 174 302 175
rect 302 174 303 175
rect 303 174 304 175
rect 304 174 305 175
rect 305 174 306 175
rect 306 174 307 175
rect 307 174 308 175
rect 308 174 309 175
rect 309 174 310 175
rect 310 174 311 175
rect 311 174 312 175
rect 312 174 313 175
rect 313 174 314 175
rect 314 174 315 175
rect 315 174 316 175
rect 316 174 317 175
rect 317 174 318 175
rect 348 174 349 175
rect 349 174 350 175
rect 350 174 351 175
rect 351 174 352 175
rect 352 174 353 175
rect 353 174 354 175
rect 354 174 355 175
rect 355 174 356 175
rect 134 173 135 174
rect 135 173 136 174
rect 136 173 137 174
rect 137 173 138 174
rect 138 173 139 174
rect 139 173 140 174
rect 140 173 141 174
rect 141 173 142 174
rect 142 173 143 174
rect 143 173 144 174
rect 290 173 291 174
rect 291 173 292 174
rect 292 173 293 174
rect 293 173 294 174
rect 294 173 295 174
rect 295 173 296 174
rect 296 173 297 174
rect 297 173 298 174
rect 298 173 299 174
rect 299 173 300 174
rect 300 173 301 174
rect 301 173 302 174
rect 302 173 303 174
rect 303 173 304 174
rect 304 173 305 174
rect 305 173 306 174
rect 306 173 307 174
rect 307 173 308 174
rect 308 173 309 174
rect 309 173 310 174
rect 310 173 311 174
rect 311 173 312 174
rect 312 173 313 174
rect 313 173 314 174
rect 314 173 315 174
rect 315 173 316 174
rect 316 173 317 174
rect 317 173 318 174
rect 348 173 349 174
rect 349 173 350 174
rect 350 173 351 174
rect 351 173 352 174
rect 352 173 353 174
rect 353 173 354 174
rect 354 173 355 174
rect 135 172 136 173
rect 136 172 137 173
rect 137 172 138 173
rect 138 172 139 173
rect 139 172 140 173
rect 140 172 141 173
rect 141 172 142 173
rect 142 172 143 173
rect 143 172 144 173
rect 144 172 145 173
rect 289 172 290 173
rect 290 172 291 173
rect 291 172 292 173
rect 292 172 293 173
rect 293 172 294 173
rect 294 172 295 173
rect 295 172 296 173
rect 296 172 297 173
rect 297 172 298 173
rect 298 172 299 173
rect 299 172 300 173
rect 300 172 301 173
rect 301 172 302 173
rect 302 172 303 173
rect 303 172 304 173
rect 304 172 305 173
rect 305 172 306 173
rect 306 172 307 173
rect 307 172 308 173
rect 308 172 309 173
rect 309 172 310 173
rect 310 172 311 173
rect 311 172 312 173
rect 312 172 313 173
rect 313 172 314 173
rect 314 172 315 173
rect 315 172 316 173
rect 316 172 317 173
rect 317 172 318 173
rect 349 172 350 173
rect 350 172 351 173
rect 351 172 352 173
rect 352 172 353 173
rect 353 172 354 173
rect 354 172 355 173
rect 135 171 136 172
rect 136 171 137 172
rect 137 171 138 172
rect 138 171 139 172
rect 139 171 140 172
rect 140 171 141 172
rect 141 171 142 172
rect 142 171 143 172
rect 143 171 144 172
rect 144 171 145 172
rect 289 171 290 172
rect 290 171 291 172
rect 291 171 292 172
rect 292 171 293 172
rect 293 171 294 172
rect 294 171 295 172
rect 295 171 296 172
rect 296 171 297 172
rect 297 171 298 172
rect 298 171 299 172
rect 299 171 300 172
rect 300 171 301 172
rect 301 171 302 172
rect 302 171 303 172
rect 303 171 304 172
rect 304 171 305 172
rect 305 171 306 172
rect 306 171 307 172
rect 307 171 308 172
rect 308 171 309 172
rect 309 171 310 172
rect 310 171 311 172
rect 312 171 313 172
rect 313 171 314 172
rect 314 171 315 172
rect 315 171 316 172
rect 316 171 317 172
rect 317 171 318 172
rect 349 171 350 172
rect 350 171 351 172
rect 351 171 352 172
rect 352 171 353 172
rect 353 171 354 172
rect 354 171 355 172
rect 136 170 137 171
rect 137 170 138 171
rect 138 170 139 171
rect 139 170 140 171
rect 140 170 141 171
rect 141 170 142 171
rect 142 170 143 171
rect 143 170 144 171
rect 144 170 145 171
rect 145 170 146 171
rect 288 170 289 171
rect 289 170 290 171
rect 290 170 291 171
rect 291 170 292 171
rect 292 170 293 171
rect 293 170 294 171
rect 294 170 295 171
rect 295 170 296 171
rect 296 170 297 171
rect 297 170 298 171
rect 298 170 299 171
rect 299 170 300 171
rect 300 170 301 171
rect 301 170 302 171
rect 302 170 303 171
rect 303 170 304 171
rect 304 170 305 171
rect 305 170 306 171
rect 306 170 307 171
rect 307 170 308 171
rect 308 170 309 171
rect 312 170 313 171
rect 313 170 314 171
rect 314 170 315 171
rect 315 170 316 171
rect 316 170 317 171
rect 317 170 318 171
rect 349 170 350 171
rect 350 170 351 171
rect 351 170 352 171
rect 352 170 353 171
rect 353 170 354 171
rect 354 170 355 171
rect 136 169 137 170
rect 137 169 138 170
rect 138 169 139 170
rect 139 169 140 170
rect 140 169 141 170
rect 141 169 142 170
rect 142 169 143 170
rect 143 169 144 170
rect 144 169 145 170
rect 145 169 146 170
rect 288 169 289 170
rect 289 169 290 170
rect 290 169 291 170
rect 291 169 292 170
rect 292 169 293 170
rect 293 169 294 170
rect 294 169 295 170
rect 295 169 296 170
rect 296 169 297 170
rect 297 169 298 170
rect 298 169 299 170
rect 299 169 300 170
rect 300 169 301 170
rect 301 169 302 170
rect 302 169 303 170
rect 303 169 304 170
rect 304 169 305 170
rect 305 169 306 170
rect 306 169 307 170
rect 312 169 313 170
rect 313 169 314 170
rect 314 169 315 170
rect 315 169 316 170
rect 316 169 317 170
rect 317 169 318 170
rect 349 169 350 170
rect 350 169 351 170
rect 351 169 352 170
rect 352 169 353 170
rect 353 169 354 170
rect 354 169 355 170
rect 137 168 138 169
rect 138 168 139 169
rect 139 168 140 169
rect 140 168 141 169
rect 141 168 142 169
rect 142 168 143 169
rect 143 168 144 169
rect 144 168 145 169
rect 145 168 146 169
rect 146 168 147 169
rect 287 168 288 169
rect 288 168 289 169
rect 289 168 290 169
rect 290 168 291 169
rect 291 168 292 169
rect 292 168 293 169
rect 293 168 294 169
rect 294 168 295 169
rect 295 168 296 169
rect 296 168 297 169
rect 297 168 298 169
rect 298 168 299 169
rect 299 168 300 169
rect 300 168 301 169
rect 301 168 302 169
rect 312 168 313 169
rect 313 168 314 169
rect 314 168 315 169
rect 315 168 316 169
rect 316 168 317 169
rect 317 168 318 169
rect 349 168 350 169
rect 350 168 351 169
rect 351 168 352 169
rect 352 168 353 169
rect 353 168 354 169
rect 354 168 355 169
rect 137 167 138 168
rect 138 167 139 168
rect 139 167 140 168
rect 140 167 141 168
rect 141 167 142 168
rect 142 167 143 168
rect 143 167 144 168
rect 144 167 145 168
rect 145 167 146 168
rect 146 167 147 168
rect 147 167 148 168
rect 286 167 287 168
rect 287 167 288 168
rect 288 167 289 168
rect 289 167 290 168
rect 290 167 291 168
rect 291 167 292 168
rect 292 167 293 168
rect 293 167 294 168
rect 294 167 295 168
rect 312 167 313 168
rect 313 167 314 168
rect 314 167 315 168
rect 315 167 316 168
rect 316 167 317 168
rect 317 167 318 168
rect 349 167 350 168
rect 350 167 351 168
rect 351 167 352 168
rect 352 167 353 168
rect 353 167 354 168
rect 354 167 355 168
rect 355 167 356 168
rect 138 166 139 167
rect 139 166 140 167
rect 140 166 141 167
rect 141 166 142 167
rect 142 166 143 167
rect 143 166 144 167
rect 144 166 145 167
rect 145 166 146 167
rect 146 166 147 167
rect 147 166 148 167
rect 286 166 287 167
rect 287 166 288 167
rect 288 166 289 167
rect 289 166 290 167
rect 290 166 291 167
rect 291 166 292 167
rect 292 166 293 167
rect 293 166 294 167
rect 294 166 295 167
rect 312 166 313 167
rect 313 166 314 167
rect 314 166 315 167
rect 315 166 316 167
rect 316 166 317 167
rect 317 166 318 167
rect 349 166 350 167
rect 350 166 351 167
rect 351 166 352 167
rect 352 166 353 167
rect 353 166 354 167
rect 354 166 355 167
rect 355 166 356 167
rect 138 165 139 166
rect 139 165 140 166
rect 140 165 141 166
rect 141 165 142 166
rect 142 165 143 166
rect 143 165 144 166
rect 144 165 145 166
rect 145 165 146 166
rect 146 165 147 166
rect 147 165 148 166
rect 148 165 149 166
rect 285 165 286 166
rect 286 165 287 166
rect 287 165 288 166
rect 288 165 289 166
rect 289 165 290 166
rect 290 165 291 166
rect 291 165 292 166
rect 292 165 293 166
rect 293 165 294 166
rect 312 165 313 166
rect 313 165 314 166
rect 314 165 315 166
rect 315 165 316 166
rect 316 165 317 166
rect 317 165 318 166
rect 349 165 350 166
rect 350 165 351 166
rect 351 165 352 166
rect 352 165 353 166
rect 353 165 354 166
rect 354 165 355 166
rect 355 165 356 166
rect 139 164 140 165
rect 140 164 141 165
rect 141 164 142 165
rect 142 164 143 165
rect 143 164 144 165
rect 144 164 145 165
rect 145 164 146 165
rect 146 164 147 165
rect 147 164 148 165
rect 148 164 149 165
rect 285 164 286 165
rect 286 164 287 165
rect 287 164 288 165
rect 288 164 289 165
rect 289 164 290 165
rect 290 164 291 165
rect 291 164 292 165
rect 292 164 293 165
rect 293 164 294 165
rect 312 164 313 165
rect 313 164 314 165
rect 314 164 315 165
rect 315 164 316 165
rect 316 164 317 165
rect 317 164 318 165
rect 349 164 350 165
rect 350 164 351 165
rect 351 164 352 165
rect 352 164 353 165
rect 353 164 354 165
rect 354 164 355 165
rect 355 164 356 165
rect 139 163 140 164
rect 140 163 141 164
rect 141 163 142 164
rect 142 163 143 164
rect 143 163 144 164
rect 144 163 145 164
rect 145 163 146 164
rect 146 163 147 164
rect 147 163 148 164
rect 148 163 149 164
rect 149 163 150 164
rect 284 163 285 164
rect 285 163 286 164
rect 286 163 287 164
rect 287 163 288 164
rect 288 163 289 164
rect 289 163 290 164
rect 290 163 291 164
rect 291 163 292 164
rect 292 163 293 164
rect 313 163 314 164
rect 314 163 315 164
rect 315 163 316 164
rect 316 163 317 164
rect 317 163 318 164
rect 349 163 350 164
rect 350 163 351 164
rect 351 163 352 164
rect 352 163 353 164
rect 353 163 354 164
rect 354 163 355 164
rect 355 163 356 164
rect 140 162 141 163
rect 141 162 142 163
rect 142 162 143 163
rect 143 162 144 163
rect 144 162 145 163
rect 145 162 146 163
rect 146 162 147 163
rect 147 162 148 163
rect 148 162 149 163
rect 149 162 150 163
rect 283 162 284 163
rect 284 162 285 163
rect 285 162 286 163
rect 286 162 287 163
rect 287 162 288 163
rect 288 162 289 163
rect 289 162 290 163
rect 290 162 291 163
rect 291 162 292 163
rect 292 162 293 163
rect 313 162 314 163
rect 314 162 315 163
rect 315 162 316 163
rect 316 162 317 163
rect 317 162 318 163
rect 318 162 319 163
rect 349 162 350 163
rect 350 162 351 163
rect 351 162 352 163
rect 352 162 353 163
rect 353 162 354 163
rect 354 162 355 163
rect 141 161 142 162
rect 142 161 143 162
rect 143 161 144 162
rect 144 161 145 162
rect 145 161 146 162
rect 146 161 147 162
rect 147 161 148 162
rect 148 161 149 162
rect 149 161 150 162
rect 150 161 151 162
rect 282 161 283 162
rect 283 161 284 162
rect 284 161 285 162
rect 285 161 286 162
rect 286 161 287 162
rect 287 161 288 162
rect 288 161 289 162
rect 289 161 290 162
rect 290 161 291 162
rect 291 161 292 162
rect 312 161 313 162
rect 313 161 314 162
rect 314 161 315 162
rect 315 161 316 162
rect 316 161 317 162
rect 317 161 318 162
rect 318 161 319 162
rect 349 161 350 162
rect 350 161 351 162
rect 351 161 352 162
rect 352 161 353 162
rect 353 161 354 162
rect 354 161 355 162
rect 141 160 142 161
rect 142 160 143 161
rect 143 160 144 161
rect 144 160 145 161
rect 145 160 146 161
rect 146 160 147 161
rect 147 160 148 161
rect 148 160 149 161
rect 149 160 150 161
rect 150 160 151 161
rect 281 160 282 161
rect 282 160 283 161
rect 283 160 284 161
rect 284 160 285 161
rect 285 160 286 161
rect 286 160 287 161
rect 287 160 288 161
rect 288 160 289 161
rect 289 160 290 161
rect 290 160 291 161
rect 312 160 313 161
rect 313 160 314 161
rect 314 160 315 161
rect 315 160 316 161
rect 316 160 317 161
rect 317 160 318 161
rect 318 160 319 161
rect 349 160 350 161
rect 350 160 351 161
rect 351 160 352 161
rect 352 160 353 161
rect 353 160 354 161
rect 354 160 355 161
rect 142 159 143 160
rect 143 159 144 160
rect 144 159 145 160
rect 145 159 146 160
rect 146 159 147 160
rect 147 159 148 160
rect 148 159 149 160
rect 149 159 150 160
rect 150 159 151 160
rect 151 159 152 160
rect 280 159 281 160
rect 281 159 282 160
rect 282 159 283 160
rect 283 159 284 160
rect 284 159 285 160
rect 285 159 286 160
rect 286 159 287 160
rect 287 159 288 160
rect 288 159 289 160
rect 289 159 290 160
rect 290 159 291 160
rect 311 159 312 160
rect 312 159 313 160
rect 313 159 314 160
rect 314 159 315 160
rect 315 159 316 160
rect 316 159 317 160
rect 317 159 318 160
rect 318 159 319 160
rect 349 159 350 160
rect 350 159 351 160
rect 351 159 352 160
rect 352 159 353 160
rect 353 159 354 160
rect 354 159 355 160
rect 355 159 356 160
rect 356 159 357 160
rect 142 158 143 159
rect 143 158 144 159
rect 144 158 145 159
rect 145 158 146 159
rect 146 158 147 159
rect 147 158 148 159
rect 148 158 149 159
rect 149 158 150 159
rect 150 158 151 159
rect 151 158 152 159
rect 279 158 280 159
rect 280 158 281 159
rect 281 158 282 159
rect 282 158 283 159
rect 283 158 284 159
rect 284 158 285 159
rect 285 158 286 159
rect 286 158 287 159
rect 287 158 288 159
rect 288 158 289 159
rect 289 158 290 159
rect 311 158 312 159
rect 312 158 313 159
rect 313 158 314 159
rect 314 158 315 159
rect 315 158 316 159
rect 316 158 317 159
rect 317 158 318 159
rect 318 158 319 159
rect 349 158 350 159
rect 350 158 351 159
rect 351 158 352 159
rect 352 158 353 159
rect 353 158 354 159
rect 354 158 355 159
rect 355 158 356 159
rect 356 158 357 159
rect 357 158 358 159
rect 358 158 359 159
rect 143 157 144 158
rect 144 157 145 158
rect 145 157 146 158
rect 146 157 147 158
rect 147 157 148 158
rect 148 157 149 158
rect 149 157 150 158
rect 150 157 151 158
rect 151 157 152 158
rect 152 157 153 158
rect 278 157 279 158
rect 279 157 280 158
rect 280 157 281 158
rect 281 157 282 158
rect 282 157 283 158
rect 283 157 284 158
rect 284 157 285 158
rect 285 157 286 158
rect 286 157 287 158
rect 287 157 288 158
rect 288 157 289 158
rect 311 157 312 158
rect 312 157 313 158
rect 313 157 314 158
rect 314 157 315 158
rect 315 157 316 158
rect 316 157 317 158
rect 317 157 318 158
rect 318 157 319 158
rect 349 157 350 158
rect 350 157 351 158
rect 351 157 352 158
rect 352 157 353 158
rect 353 157 354 158
rect 354 157 355 158
rect 355 157 356 158
rect 356 157 357 158
rect 357 157 358 158
rect 358 157 359 158
rect 143 156 144 157
rect 144 156 145 157
rect 145 156 146 157
rect 146 156 147 157
rect 147 156 148 157
rect 148 156 149 157
rect 149 156 150 157
rect 150 156 151 157
rect 151 156 152 157
rect 152 156 153 157
rect 277 156 278 157
rect 278 156 279 157
rect 279 156 280 157
rect 280 156 281 157
rect 281 156 282 157
rect 282 156 283 157
rect 283 156 284 157
rect 284 156 285 157
rect 285 156 286 157
rect 286 156 287 157
rect 287 156 288 157
rect 310 156 311 157
rect 311 156 312 157
rect 312 156 313 157
rect 313 156 314 157
rect 314 156 315 157
rect 315 156 316 157
rect 316 156 317 157
rect 317 156 318 157
rect 318 156 319 157
rect 319 156 320 157
rect 349 156 350 157
rect 350 156 351 157
rect 351 156 352 157
rect 352 156 353 157
rect 353 156 354 157
rect 354 156 355 157
rect 355 156 356 157
rect 356 156 357 157
rect 357 156 358 157
rect 358 156 359 157
rect 359 156 360 157
rect 144 155 145 156
rect 145 155 146 156
rect 146 155 147 156
rect 147 155 148 156
rect 148 155 149 156
rect 149 155 150 156
rect 150 155 151 156
rect 151 155 152 156
rect 152 155 153 156
rect 153 155 154 156
rect 275 155 276 156
rect 276 155 277 156
rect 277 155 278 156
rect 278 155 279 156
rect 279 155 280 156
rect 280 155 281 156
rect 281 155 282 156
rect 282 155 283 156
rect 283 155 284 156
rect 284 155 285 156
rect 285 155 286 156
rect 286 155 287 156
rect 287 155 288 156
rect 310 155 311 156
rect 311 155 312 156
rect 312 155 313 156
rect 313 155 314 156
rect 314 155 315 156
rect 315 155 316 156
rect 316 155 317 156
rect 317 155 318 156
rect 318 155 319 156
rect 319 155 320 156
rect 349 155 350 156
rect 350 155 351 156
rect 351 155 352 156
rect 352 155 353 156
rect 353 155 354 156
rect 354 155 355 156
rect 355 155 356 156
rect 356 155 357 156
rect 357 155 358 156
rect 358 155 359 156
rect 359 155 360 156
rect 144 154 145 155
rect 145 154 146 155
rect 146 154 147 155
rect 147 154 148 155
rect 148 154 149 155
rect 149 154 150 155
rect 150 154 151 155
rect 151 154 152 155
rect 152 154 153 155
rect 153 154 154 155
rect 154 154 155 155
rect 274 154 275 155
rect 275 154 276 155
rect 276 154 277 155
rect 277 154 278 155
rect 278 154 279 155
rect 279 154 280 155
rect 280 154 281 155
rect 281 154 282 155
rect 282 154 283 155
rect 283 154 284 155
rect 284 154 285 155
rect 285 154 286 155
rect 286 154 287 155
rect 309 154 310 155
rect 310 154 311 155
rect 311 154 312 155
rect 312 154 313 155
rect 313 154 314 155
rect 314 154 315 155
rect 315 154 316 155
rect 316 154 317 155
rect 317 154 318 155
rect 318 154 319 155
rect 319 154 320 155
rect 349 154 350 155
rect 350 154 351 155
rect 351 154 352 155
rect 352 154 353 155
rect 353 154 354 155
rect 354 154 355 155
rect 355 154 356 155
rect 356 154 357 155
rect 357 154 358 155
rect 358 154 359 155
rect 359 154 360 155
rect 360 154 361 155
rect 145 153 146 154
rect 146 153 147 154
rect 147 153 148 154
rect 148 153 149 154
rect 149 153 150 154
rect 150 153 151 154
rect 151 153 152 154
rect 152 153 153 154
rect 153 153 154 154
rect 154 153 155 154
rect 155 153 156 154
rect 273 153 274 154
rect 274 153 275 154
rect 275 153 276 154
rect 276 153 277 154
rect 277 153 278 154
rect 278 153 279 154
rect 279 153 280 154
rect 280 153 281 154
rect 281 153 282 154
rect 282 153 283 154
rect 283 153 284 154
rect 284 153 285 154
rect 285 153 286 154
rect 308 153 309 154
rect 309 153 310 154
rect 310 153 311 154
rect 311 153 312 154
rect 312 153 313 154
rect 313 153 314 154
rect 314 153 315 154
rect 315 153 316 154
rect 316 153 317 154
rect 317 153 318 154
rect 318 153 319 154
rect 319 153 320 154
rect 320 153 321 154
rect 348 153 349 154
rect 349 153 350 154
rect 350 153 351 154
rect 351 153 352 154
rect 352 153 353 154
rect 353 153 354 154
rect 354 153 355 154
rect 355 153 356 154
rect 356 153 357 154
rect 357 153 358 154
rect 358 153 359 154
rect 359 153 360 154
rect 360 153 361 154
rect 146 152 147 153
rect 147 152 148 153
rect 148 152 149 153
rect 149 152 150 153
rect 150 152 151 153
rect 151 152 152 153
rect 152 152 153 153
rect 153 152 154 153
rect 154 152 155 153
rect 155 152 156 153
rect 156 152 157 153
rect 157 152 158 153
rect 272 152 273 153
rect 273 152 274 153
rect 274 152 275 153
rect 275 152 276 153
rect 276 152 277 153
rect 277 152 278 153
rect 278 152 279 153
rect 279 152 280 153
rect 280 152 281 153
rect 281 152 282 153
rect 282 152 283 153
rect 283 152 284 153
rect 284 152 285 153
rect 308 152 309 153
rect 309 152 310 153
rect 310 152 311 153
rect 311 152 312 153
rect 312 152 313 153
rect 313 152 314 153
rect 314 152 315 153
rect 315 152 316 153
rect 316 152 317 153
rect 317 152 318 153
rect 318 152 319 153
rect 319 152 320 153
rect 320 152 321 153
rect 348 152 349 153
rect 349 152 350 153
rect 350 152 351 153
rect 354 152 355 153
rect 355 152 356 153
rect 356 152 357 153
rect 357 152 358 153
rect 358 152 359 153
rect 359 152 360 153
rect 360 152 361 153
rect 146 151 147 152
rect 147 151 148 152
rect 148 151 149 152
rect 149 151 150 152
rect 150 151 151 152
rect 151 151 152 152
rect 152 151 153 152
rect 153 151 154 152
rect 154 151 155 152
rect 155 151 156 152
rect 156 151 157 152
rect 157 151 158 152
rect 158 151 159 152
rect 159 151 160 152
rect 175 151 176 152
rect 176 151 177 152
rect 177 151 178 152
rect 178 151 179 152
rect 270 151 271 152
rect 271 151 272 152
rect 272 151 273 152
rect 273 151 274 152
rect 274 151 275 152
rect 275 151 276 152
rect 276 151 277 152
rect 277 151 278 152
rect 278 151 279 152
rect 279 151 280 152
rect 280 151 281 152
rect 281 151 282 152
rect 282 151 283 152
rect 283 151 284 152
rect 307 151 308 152
rect 308 151 309 152
rect 309 151 310 152
rect 310 151 311 152
rect 311 151 312 152
rect 312 151 313 152
rect 313 151 314 152
rect 314 151 315 152
rect 315 151 316 152
rect 316 151 317 152
rect 317 151 318 152
rect 318 151 319 152
rect 319 151 320 152
rect 320 151 321 152
rect 348 151 349 152
rect 349 151 350 152
rect 350 151 351 152
rect 355 151 356 152
rect 356 151 357 152
rect 357 151 358 152
rect 358 151 359 152
rect 359 151 360 152
rect 360 151 361 152
rect 361 151 362 152
rect 362 151 363 152
rect 363 151 364 152
rect 147 150 148 151
rect 148 150 149 151
rect 149 150 150 151
rect 150 150 151 151
rect 151 150 152 151
rect 152 150 153 151
rect 153 150 154 151
rect 154 150 155 151
rect 155 150 156 151
rect 156 150 157 151
rect 157 150 158 151
rect 158 150 159 151
rect 159 150 160 151
rect 160 150 161 151
rect 161 150 162 151
rect 162 150 163 151
rect 163 150 164 151
rect 164 150 165 151
rect 165 150 166 151
rect 166 150 167 151
rect 167 150 168 151
rect 168 150 169 151
rect 169 150 170 151
rect 170 150 171 151
rect 171 150 172 151
rect 172 150 173 151
rect 173 150 174 151
rect 174 150 175 151
rect 175 150 176 151
rect 176 150 177 151
rect 177 150 178 151
rect 178 150 179 151
rect 269 150 270 151
rect 270 150 271 151
rect 271 150 272 151
rect 272 150 273 151
rect 273 150 274 151
rect 274 150 275 151
rect 275 150 276 151
rect 276 150 277 151
rect 277 150 278 151
rect 278 150 279 151
rect 279 150 280 151
rect 280 150 281 151
rect 281 150 282 151
rect 282 150 283 151
rect 307 150 308 151
rect 308 150 309 151
rect 309 150 310 151
rect 310 150 311 151
rect 311 150 312 151
rect 312 150 313 151
rect 313 150 314 151
rect 314 150 315 151
rect 315 150 316 151
rect 316 150 317 151
rect 317 150 318 151
rect 318 150 319 151
rect 319 150 320 151
rect 320 150 321 151
rect 321 150 322 151
rect 348 150 349 151
rect 349 150 350 151
rect 356 150 357 151
rect 357 150 358 151
rect 358 150 359 151
rect 359 150 360 151
rect 360 150 361 151
rect 361 150 362 151
rect 362 150 363 151
rect 363 150 364 151
rect 364 150 365 151
rect 148 149 149 150
rect 149 149 150 150
rect 150 149 151 150
rect 151 149 152 150
rect 152 149 153 150
rect 153 149 154 150
rect 154 149 155 150
rect 155 149 156 150
rect 156 149 157 150
rect 157 149 158 150
rect 158 149 159 150
rect 159 149 160 150
rect 160 149 161 150
rect 161 149 162 150
rect 162 149 163 150
rect 163 149 164 150
rect 164 149 165 150
rect 165 149 166 150
rect 166 149 167 150
rect 167 149 168 150
rect 168 149 169 150
rect 169 149 170 150
rect 170 149 171 150
rect 171 149 172 150
rect 172 149 173 150
rect 173 149 174 150
rect 174 149 175 150
rect 175 149 176 150
rect 176 149 177 150
rect 177 149 178 150
rect 178 149 179 150
rect 179 149 180 150
rect 268 149 269 150
rect 269 149 270 150
rect 270 149 271 150
rect 271 149 272 150
rect 272 149 273 150
rect 273 149 274 150
rect 274 149 275 150
rect 275 149 276 150
rect 276 149 277 150
rect 277 149 278 150
rect 278 149 279 150
rect 279 149 280 150
rect 280 149 281 150
rect 306 149 307 150
rect 307 149 308 150
rect 308 149 309 150
rect 309 149 310 150
rect 310 149 311 150
rect 311 149 312 150
rect 312 149 313 150
rect 313 149 314 150
rect 315 149 316 150
rect 316 149 317 150
rect 317 149 318 150
rect 318 149 319 150
rect 319 149 320 150
rect 320 149 321 150
rect 321 149 322 150
rect 347 149 348 150
rect 348 149 349 150
rect 349 149 350 150
rect 356 149 357 150
rect 357 149 358 150
rect 358 149 359 150
rect 359 149 360 150
rect 360 149 361 150
rect 361 149 362 150
rect 362 149 363 150
rect 363 149 364 150
rect 364 149 365 150
rect 365 149 366 150
rect 366 149 367 150
rect 149 148 150 149
rect 150 148 151 149
rect 151 148 152 149
rect 152 148 153 149
rect 153 148 154 149
rect 154 148 155 149
rect 155 148 156 149
rect 156 148 157 149
rect 157 148 158 149
rect 158 148 159 149
rect 159 148 160 149
rect 160 148 161 149
rect 161 148 162 149
rect 162 148 163 149
rect 163 148 164 149
rect 164 148 165 149
rect 165 148 166 149
rect 166 148 167 149
rect 167 148 168 149
rect 168 148 169 149
rect 169 148 170 149
rect 170 148 171 149
rect 171 148 172 149
rect 172 148 173 149
rect 173 148 174 149
rect 174 148 175 149
rect 175 148 176 149
rect 176 148 177 149
rect 177 148 178 149
rect 178 148 179 149
rect 179 148 180 149
rect 180 148 181 149
rect 181 148 182 149
rect 266 148 267 149
rect 267 148 268 149
rect 268 148 269 149
rect 269 148 270 149
rect 270 148 271 149
rect 271 148 272 149
rect 272 148 273 149
rect 273 148 274 149
rect 274 148 275 149
rect 275 148 276 149
rect 276 148 277 149
rect 277 148 278 149
rect 278 148 279 149
rect 279 148 280 149
rect 305 148 306 149
rect 306 148 307 149
rect 307 148 308 149
rect 308 148 309 149
rect 309 148 310 149
rect 310 148 311 149
rect 311 148 312 149
rect 312 148 313 149
rect 313 148 314 149
rect 315 148 316 149
rect 316 148 317 149
rect 317 148 318 149
rect 318 148 319 149
rect 319 148 320 149
rect 320 148 321 149
rect 321 148 322 149
rect 322 148 323 149
rect 356 148 357 149
rect 357 148 358 149
rect 358 148 359 149
rect 359 148 360 149
rect 360 148 361 149
rect 361 148 362 149
rect 362 148 363 149
rect 363 148 364 149
rect 364 148 365 149
rect 365 148 366 149
rect 366 148 367 149
rect 367 148 368 149
rect 150 147 151 148
rect 151 147 152 148
rect 152 147 153 148
rect 153 147 154 148
rect 154 147 155 148
rect 155 147 156 148
rect 156 147 157 148
rect 157 147 158 148
rect 158 147 159 148
rect 159 147 160 148
rect 160 147 161 148
rect 161 147 162 148
rect 162 147 163 148
rect 163 147 164 148
rect 164 147 165 148
rect 165 147 166 148
rect 166 147 167 148
rect 167 147 168 148
rect 168 147 169 148
rect 169 147 170 148
rect 170 147 171 148
rect 171 147 172 148
rect 172 147 173 148
rect 173 147 174 148
rect 174 147 175 148
rect 175 147 176 148
rect 176 147 177 148
rect 177 147 178 148
rect 178 147 179 148
rect 179 147 180 148
rect 180 147 181 148
rect 181 147 182 148
rect 182 147 183 148
rect 265 147 266 148
rect 266 147 267 148
rect 267 147 268 148
rect 268 147 269 148
rect 269 147 270 148
rect 270 147 271 148
rect 271 147 272 148
rect 272 147 273 148
rect 273 147 274 148
rect 274 147 275 148
rect 275 147 276 148
rect 276 147 277 148
rect 277 147 278 148
rect 278 147 279 148
rect 305 147 306 148
rect 306 147 307 148
rect 307 147 308 148
rect 308 147 309 148
rect 309 147 310 148
rect 310 147 311 148
rect 311 147 312 148
rect 312 147 313 148
rect 313 147 314 148
rect 315 147 316 148
rect 316 147 317 148
rect 317 147 318 148
rect 318 147 319 148
rect 319 147 320 148
rect 320 147 321 148
rect 321 147 322 148
rect 322 147 323 148
rect 356 147 357 148
rect 357 147 358 148
rect 358 147 359 148
rect 359 147 360 148
rect 360 147 361 148
rect 361 147 362 148
rect 362 147 363 148
rect 363 147 364 148
rect 364 147 365 148
rect 365 147 366 148
rect 366 147 367 148
rect 367 147 368 148
rect 368 147 369 148
rect 369 147 370 148
rect 152 146 153 147
rect 153 146 154 147
rect 154 146 155 147
rect 155 146 156 147
rect 156 146 157 147
rect 157 146 158 147
rect 158 146 159 147
rect 159 146 160 147
rect 160 146 161 147
rect 161 146 162 147
rect 162 146 163 147
rect 163 146 164 147
rect 164 146 165 147
rect 165 146 166 147
rect 166 146 167 147
rect 167 146 168 147
rect 168 146 169 147
rect 169 146 170 147
rect 170 146 171 147
rect 171 146 172 147
rect 172 146 173 147
rect 173 146 174 147
rect 174 146 175 147
rect 175 146 176 147
rect 176 146 177 147
rect 177 146 178 147
rect 178 146 179 147
rect 179 146 180 147
rect 180 146 181 147
rect 181 146 182 147
rect 182 146 183 147
rect 183 146 184 147
rect 263 146 264 147
rect 264 146 265 147
rect 265 146 266 147
rect 266 146 267 147
rect 267 146 268 147
rect 268 146 269 147
rect 269 146 270 147
rect 270 146 271 147
rect 271 146 272 147
rect 272 146 273 147
rect 273 146 274 147
rect 274 146 275 147
rect 275 146 276 147
rect 276 146 277 147
rect 277 146 278 147
rect 304 146 305 147
rect 305 146 306 147
rect 306 146 307 147
rect 307 146 308 147
rect 308 146 309 147
rect 309 146 310 147
rect 310 146 311 147
rect 311 146 312 147
rect 312 146 313 147
rect 316 146 317 147
rect 317 146 318 147
rect 318 146 319 147
rect 319 146 320 147
rect 320 146 321 147
rect 321 146 322 147
rect 322 146 323 147
rect 323 146 324 147
rect 356 146 357 147
rect 357 146 358 147
rect 358 146 359 147
rect 360 146 361 147
rect 361 146 362 147
rect 362 146 363 147
rect 363 146 364 147
rect 364 146 365 147
rect 365 146 366 147
rect 366 146 367 147
rect 367 146 368 147
rect 368 146 369 147
rect 369 146 370 147
rect 370 146 371 147
rect 154 145 155 146
rect 155 145 156 146
rect 156 145 157 146
rect 157 145 158 146
rect 158 145 159 146
rect 159 145 160 146
rect 160 145 161 146
rect 161 145 162 146
rect 162 145 163 146
rect 163 145 164 146
rect 164 145 165 146
rect 165 145 166 146
rect 166 145 167 146
rect 167 145 168 146
rect 168 145 169 146
rect 169 145 170 146
rect 170 145 171 146
rect 171 145 172 146
rect 172 145 173 146
rect 173 145 174 146
rect 174 145 175 146
rect 175 145 176 146
rect 176 145 177 146
rect 177 145 178 146
rect 178 145 179 146
rect 179 145 180 146
rect 180 145 181 146
rect 181 145 182 146
rect 182 145 183 146
rect 183 145 184 146
rect 184 145 185 146
rect 185 145 186 146
rect 262 145 263 146
rect 263 145 264 146
rect 264 145 265 146
rect 265 145 266 146
rect 266 145 267 146
rect 267 145 268 146
rect 268 145 269 146
rect 269 145 270 146
rect 270 145 271 146
rect 271 145 272 146
rect 272 145 273 146
rect 273 145 274 146
rect 274 145 275 146
rect 275 145 276 146
rect 276 145 277 146
rect 303 145 304 146
rect 304 145 305 146
rect 305 145 306 146
rect 306 145 307 146
rect 307 145 308 146
rect 308 145 309 146
rect 309 145 310 146
rect 310 145 311 146
rect 311 145 312 146
rect 312 145 313 146
rect 316 145 317 146
rect 317 145 318 146
rect 318 145 319 146
rect 319 145 320 146
rect 320 145 321 146
rect 321 145 322 146
rect 322 145 323 146
rect 323 145 324 146
rect 324 145 325 146
rect 356 145 357 146
rect 357 145 358 146
rect 358 145 359 146
rect 362 145 363 146
rect 363 145 364 146
rect 364 145 365 146
rect 365 145 366 146
rect 366 145 367 146
rect 367 145 368 146
rect 368 145 369 146
rect 369 145 370 146
rect 370 145 371 146
rect 371 145 372 146
rect 156 144 157 145
rect 157 144 158 145
rect 158 144 159 145
rect 159 144 160 145
rect 160 144 161 145
rect 161 144 162 145
rect 162 144 163 145
rect 163 144 164 145
rect 164 144 165 145
rect 165 144 166 145
rect 166 144 167 145
rect 167 144 168 145
rect 168 144 169 145
rect 169 144 170 145
rect 170 144 171 145
rect 171 144 172 145
rect 172 144 173 145
rect 173 144 174 145
rect 174 144 175 145
rect 175 144 176 145
rect 176 144 177 145
rect 177 144 178 145
rect 178 144 179 145
rect 179 144 180 145
rect 180 144 181 145
rect 181 144 182 145
rect 182 144 183 145
rect 183 144 184 145
rect 184 144 185 145
rect 185 144 186 145
rect 186 144 187 145
rect 187 144 188 145
rect 260 144 261 145
rect 261 144 262 145
rect 262 144 263 145
rect 263 144 264 145
rect 264 144 265 145
rect 265 144 266 145
rect 266 144 267 145
rect 267 144 268 145
rect 268 144 269 145
rect 269 144 270 145
rect 270 144 271 145
rect 271 144 272 145
rect 272 144 273 145
rect 273 144 274 145
rect 274 144 275 145
rect 303 144 304 145
rect 304 144 305 145
rect 305 144 306 145
rect 306 144 307 145
rect 307 144 308 145
rect 308 144 309 145
rect 309 144 310 145
rect 310 144 311 145
rect 311 144 312 145
rect 312 144 313 145
rect 316 144 317 145
rect 317 144 318 145
rect 318 144 319 145
rect 319 144 320 145
rect 320 144 321 145
rect 321 144 322 145
rect 322 144 323 145
rect 323 144 324 145
rect 324 144 325 145
rect 325 144 326 145
rect 364 144 365 145
rect 365 144 366 145
rect 366 144 367 145
rect 367 144 368 145
rect 368 144 369 145
rect 369 144 370 145
rect 370 144 371 145
rect 371 144 372 145
rect 372 144 373 145
rect 159 143 160 144
rect 160 143 161 144
rect 161 143 162 144
rect 162 143 163 144
rect 163 143 164 144
rect 164 143 165 144
rect 165 143 166 144
rect 166 143 167 144
rect 167 143 168 144
rect 168 143 169 144
rect 169 143 170 144
rect 170 143 171 144
rect 171 143 172 144
rect 172 143 173 144
rect 173 143 174 144
rect 174 143 175 144
rect 175 143 176 144
rect 176 143 177 144
rect 177 143 178 144
rect 178 143 179 144
rect 179 143 180 144
rect 180 143 181 144
rect 181 143 182 144
rect 182 143 183 144
rect 183 143 184 144
rect 184 143 185 144
rect 185 143 186 144
rect 186 143 187 144
rect 187 143 188 144
rect 188 143 189 144
rect 189 143 190 144
rect 190 143 191 144
rect 258 143 259 144
rect 259 143 260 144
rect 260 143 261 144
rect 261 143 262 144
rect 262 143 263 144
rect 263 143 264 144
rect 264 143 265 144
rect 265 143 266 144
rect 266 143 267 144
rect 267 143 268 144
rect 268 143 269 144
rect 269 143 270 144
rect 270 143 271 144
rect 271 143 272 144
rect 272 143 273 144
rect 273 143 274 144
rect 302 143 303 144
rect 303 143 304 144
rect 304 143 305 144
rect 305 143 306 144
rect 307 143 308 144
rect 308 143 309 144
rect 309 143 310 144
rect 310 143 311 144
rect 311 143 312 144
rect 312 143 313 144
rect 313 143 314 144
rect 317 143 318 144
rect 318 143 319 144
rect 319 143 320 144
rect 320 143 321 144
rect 321 143 322 144
rect 322 143 323 144
rect 323 143 324 144
rect 324 143 325 144
rect 325 143 326 144
rect 326 143 327 144
rect 365 143 366 144
rect 366 143 367 144
rect 367 143 368 144
rect 368 143 369 144
rect 369 143 370 144
rect 370 143 371 144
rect 371 143 372 144
rect 372 143 373 144
rect 373 143 374 144
rect 162 142 163 143
rect 163 142 164 143
rect 164 142 165 143
rect 165 142 166 143
rect 166 142 167 143
rect 167 142 168 143
rect 168 142 169 143
rect 169 142 170 143
rect 170 142 171 143
rect 171 142 172 143
rect 172 142 173 143
rect 173 142 174 143
rect 174 142 175 143
rect 175 142 176 143
rect 176 142 177 143
rect 177 142 178 143
rect 178 142 179 143
rect 179 142 180 143
rect 180 142 181 143
rect 181 142 182 143
rect 182 142 183 143
rect 183 142 184 143
rect 184 142 185 143
rect 185 142 186 143
rect 186 142 187 143
rect 187 142 188 143
rect 188 142 189 143
rect 189 142 190 143
rect 190 142 191 143
rect 191 142 192 143
rect 192 142 193 143
rect 193 142 194 143
rect 194 142 195 143
rect 256 142 257 143
rect 257 142 258 143
rect 258 142 259 143
rect 259 142 260 143
rect 260 142 261 143
rect 261 142 262 143
rect 262 142 263 143
rect 263 142 264 143
rect 264 142 265 143
rect 265 142 266 143
rect 266 142 267 143
rect 267 142 268 143
rect 268 142 269 143
rect 269 142 270 143
rect 270 142 271 143
rect 271 142 272 143
rect 272 142 273 143
rect 301 142 302 143
rect 302 142 303 143
rect 303 142 304 143
rect 304 142 305 143
rect 307 142 308 143
rect 308 142 309 143
rect 309 142 310 143
rect 310 142 311 143
rect 311 142 312 143
rect 312 142 313 143
rect 313 142 314 143
rect 317 142 318 143
rect 318 142 319 143
rect 319 142 320 143
rect 320 142 321 143
rect 321 142 322 143
rect 322 142 323 143
rect 323 142 324 143
rect 324 142 325 143
rect 325 142 326 143
rect 326 142 327 143
rect 327 142 328 143
rect 367 142 368 143
rect 368 142 369 143
rect 369 142 370 143
rect 370 142 371 143
rect 371 142 372 143
rect 372 142 373 143
rect 373 142 374 143
rect 374 142 375 143
rect 179 141 180 142
rect 180 141 181 142
rect 181 141 182 142
rect 182 141 183 142
rect 183 141 184 142
rect 184 141 185 142
rect 185 141 186 142
rect 186 141 187 142
rect 187 141 188 142
rect 188 141 189 142
rect 189 141 190 142
rect 190 141 191 142
rect 191 141 192 142
rect 192 141 193 142
rect 193 141 194 142
rect 194 141 195 142
rect 195 141 196 142
rect 196 141 197 142
rect 197 141 198 142
rect 198 141 199 142
rect 254 141 255 142
rect 255 141 256 142
rect 256 141 257 142
rect 257 141 258 142
rect 258 141 259 142
rect 259 141 260 142
rect 260 141 261 142
rect 261 141 262 142
rect 262 141 263 142
rect 263 141 264 142
rect 264 141 265 142
rect 265 141 266 142
rect 266 141 267 142
rect 267 141 268 142
rect 268 141 269 142
rect 269 141 270 142
rect 270 141 271 142
rect 300 141 301 142
rect 301 141 302 142
rect 302 141 303 142
rect 303 141 304 142
rect 304 141 305 142
rect 307 141 308 142
rect 308 141 309 142
rect 309 141 310 142
rect 310 141 311 142
rect 311 141 312 142
rect 312 141 313 142
rect 313 141 314 142
rect 318 141 319 142
rect 319 141 320 142
rect 320 141 321 142
rect 321 141 322 142
rect 322 141 323 142
rect 323 141 324 142
rect 324 141 325 142
rect 325 141 326 142
rect 326 141 327 142
rect 327 141 328 142
rect 328 141 329 142
rect 329 141 330 142
rect 368 141 369 142
rect 369 141 370 142
rect 370 141 371 142
rect 371 141 372 142
rect 372 141 373 142
rect 373 141 374 142
rect 374 141 375 142
rect 375 141 376 142
rect 179 140 180 141
rect 180 140 181 141
rect 181 140 182 141
rect 182 140 183 141
rect 183 140 184 141
rect 184 140 185 141
rect 185 140 186 141
rect 186 140 187 141
rect 187 140 188 141
rect 188 140 189 141
rect 189 140 190 141
rect 190 140 191 141
rect 191 140 192 141
rect 192 140 193 141
rect 193 140 194 141
rect 194 140 195 141
rect 195 140 196 141
rect 196 140 197 141
rect 197 140 198 141
rect 198 140 199 141
rect 199 140 200 141
rect 200 140 201 141
rect 201 140 202 141
rect 202 140 203 141
rect 252 140 253 141
rect 253 140 254 141
rect 254 140 255 141
rect 255 140 256 141
rect 256 140 257 141
rect 257 140 258 141
rect 258 140 259 141
rect 259 140 260 141
rect 260 140 261 141
rect 261 140 262 141
rect 262 140 263 141
rect 263 140 264 141
rect 264 140 265 141
rect 265 140 266 141
rect 266 140 267 141
rect 267 140 268 141
rect 268 140 269 141
rect 269 140 270 141
rect 300 140 301 141
rect 301 140 302 141
rect 302 140 303 141
rect 303 140 304 141
rect 307 140 308 141
rect 308 140 309 141
rect 309 140 310 141
rect 310 140 311 141
rect 311 140 312 141
rect 312 140 313 141
rect 313 140 314 141
rect 318 140 319 141
rect 319 140 320 141
rect 320 140 321 141
rect 321 140 322 141
rect 322 140 323 141
rect 323 140 324 141
rect 324 140 325 141
rect 325 140 326 141
rect 326 140 327 141
rect 327 140 328 141
rect 328 140 329 141
rect 329 140 330 141
rect 330 140 331 141
rect 331 140 332 141
rect 368 140 369 141
rect 369 140 370 141
rect 370 140 371 141
rect 371 140 372 141
rect 372 140 373 141
rect 373 140 374 141
rect 374 140 375 141
rect 375 140 376 141
rect 180 139 181 140
rect 181 139 182 140
rect 182 139 183 140
rect 183 139 184 140
rect 184 139 185 140
rect 185 139 186 140
rect 186 139 187 140
rect 187 139 188 140
rect 188 139 189 140
rect 189 139 190 140
rect 190 139 191 140
rect 191 139 192 140
rect 192 139 193 140
rect 193 139 194 140
rect 194 139 195 140
rect 195 139 196 140
rect 196 139 197 140
rect 197 139 198 140
rect 198 139 199 140
rect 199 139 200 140
rect 200 139 201 140
rect 201 139 202 140
rect 202 139 203 140
rect 203 139 204 140
rect 204 139 205 140
rect 205 139 206 140
rect 206 139 207 140
rect 207 139 208 140
rect 250 139 251 140
rect 251 139 252 140
rect 252 139 253 140
rect 253 139 254 140
rect 254 139 255 140
rect 255 139 256 140
rect 256 139 257 140
rect 257 139 258 140
rect 258 139 259 140
rect 259 139 260 140
rect 260 139 261 140
rect 261 139 262 140
rect 262 139 263 140
rect 263 139 264 140
rect 264 139 265 140
rect 265 139 266 140
rect 266 139 267 140
rect 267 139 268 140
rect 268 139 269 140
rect 299 139 300 140
rect 300 139 301 140
rect 301 139 302 140
rect 302 139 303 140
rect 303 139 304 140
rect 307 139 308 140
rect 308 139 309 140
rect 309 139 310 140
rect 310 139 311 140
rect 311 139 312 140
rect 312 139 313 140
rect 313 139 314 140
rect 319 139 320 140
rect 320 139 321 140
rect 321 139 322 140
rect 322 139 323 140
rect 323 139 324 140
rect 324 139 325 140
rect 325 139 326 140
rect 326 139 327 140
rect 327 139 328 140
rect 328 139 329 140
rect 329 139 330 140
rect 330 139 331 140
rect 331 139 332 140
rect 332 139 333 140
rect 333 139 334 140
rect 334 139 335 140
rect 335 139 336 140
rect 336 139 337 140
rect 369 139 370 140
rect 370 139 371 140
rect 371 139 372 140
rect 372 139 373 140
rect 373 139 374 140
rect 374 139 375 140
rect 375 139 376 140
rect 376 139 377 140
rect 180 138 181 139
rect 181 138 182 139
rect 182 138 183 139
rect 183 138 184 139
rect 184 138 185 139
rect 185 138 186 139
rect 186 138 187 139
rect 187 138 188 139
rect 188 138 189 139
rect 189 138 190 139
rect 190 138 191 139
rect 191 138 192 139
rect 192 138 193 139
rect 193 138 194 139
rect 194 138 195 139
rect 195 138 196 139
rect 196 138 197 139
rect 197 138 198 139
rect 198 138 199 139
rect 199 138 200 139
rect 200 138 201 139
rect 201 138 202 139
rect 202 138 203 139
rect 203 138 204 139
rect 204 138 205 139
rect 205 138 206 139
rect 206 138 207 139
rect 207 138 208 139
rect 208 138 209 139
rect 209 138 210 139
rect 210 138 211 139
rect 211 138 212 139
rect 247 138 248 139
rect 248 138 249 139
rect 249 138 250 139
rect 250 138 251 139
rect 251 138 252 139
rect 252 138 253 139
rect 253 138 254 139
rect 254 138 255 139
rect 255 138 256 139
rect 256 138 257 139
rect 257 138 258 139
rect 258 138 259 139
rect 259 138 260 139
rect 260 138 261 139
rect 261 138 262 139
rect 262 138 263 139
rect 263 138 264 139
rect 264 138 265 139
rect 265 138 266 139
rect 266 138 267 139
rect 298 138 299 139
rect 299 138 300 139
rect 300 138 301 139
rect 301 138 302 139
rect 302 138 303 139
rect 307 138 308 139
rect 308 138 309 139
rect 309 138 310 139
rect 310 138 311 139
rect 311 138 312 139
rect 312 138 313 139
rect 313 138 314 139
rect 320 138 321 139
rect 321 138 322 139
rect 322 138 323 139
rect 323 138 324 139
rect 324 138 325 139
rect 325 138 326 139
rect 326 138 327 139
rect 327 138 328 139
rect 328 138 329 139
rect 329 138 330 139
rect 330 138 331 139
rect 331 138 332 139
rect 332 138 333 139
rect 333 138 334 139
rect 334 138 335 139
rect 335 138 336 139
rect 336 138 337 139
rect 337 138 338 139
rect 338 138 339 139
rect 339 138 340 139
rect 340 138 341 139
rect 341 138 342 139
rect 370 138 371 139
rect 371 138 372 139
rect 372 138 373 139
rect 373 138 374 139
rect 374 138 375 139
rect 375 138 376 139
rect 376 138 377 139
rect 181 137 182 138
rect 182 137 183 138
rect 183 137 184 138
rect 184 137 185 138
rect 185 137 186 138
rect 186 137 187 138
rect 187 137 188 138
rect 188 137 189 138
rect 189 137 190 138
rect 190 137 191 138
rect 191 137 192 138
rect 192 137 193 138
rect 193 137 194 138
rect 194 137 195 138
rect 195 137 196 138
rect 196 137 197 138
rect 197 137 198 138
rect 198 137 199 138
rect 199 137 200 138
rect 200 137 201 138
rect 201 137 202 138
rect 202 137 203 138
rect 203 137 204 138
rect 204 137 205 138
rect 205 137 206 138
rect 206 137 207 138
rect 207 137 208 138
rect 208 137 209 138
rect 209 137 210 138
rect 210 137 211 138
rect 211 137 212 138
rect 212 137 213 138
rect 213 137 214 138
rect 214 137 215 138
rect 215 137 216 138
rect 244 137 245 138
rect 245 137 246 138
rect 246 137 247 138
rect 247 137 248 138
rect 248 137 249 138
rect 249 137 250 138
rect 250 137 251 138
rect 251 137 252 138
rect 252 137 253 138
rect 253 137 254 138
rect 254 137 255 138
rect 255 137 256 138
rect 256 137 257 138
rect 257 137 258 138
rect 258 137 259 138
rect 259 137 260 138
rect 260 137 261 138
rect 261 137 262 138
rect 262 137 263 138
rect 263 137 264 138
rect 264 137 265 138
rect 265 137 266 138
rect 297 137 298 138
rect 298 137 299 138
rect 299 137 300 138
rect 300 137 301 138
rect 301 137 302 138
rect 307 137 308 138
rect 308 137 309 138
rect 309 137 310 138
rect 310 137 311 138
rect 311 137 312 138
rect 312 137 313 138
rect 313 137 314 138
rect 321 137 322 138
rect 322 137 323 138
rect 323 137 324 138
rect 324 137 325 138
rect 325 137 326 138
rect 326 137 327 138
rect 327 137 328 138
rect 328 137 329 138
rect 329 137 330 138
rect 330 137 331 138
rect 331 137 332 138
rect 332 137 333 138
rect 333 137 334 138
rect 334 137 335 138
rect 335 137 336 138
rect 336 137 337 138
rect 337 137 338 138
rect 338 137 339 138
rect 339 137 340 138
rect 340 137 341 138
rect 341 137 342 138
rect 342 137 343 138
rect 343 137 344 138
rect 344 137 345 138
rect 370 137 371 138
rect 371 137 372 138
rect 372 137 373 138
rect 373 137 374 138
rect 374 137 375 138
rect 375 137 376 138
rect 376 137 377 138
rect 182 136 183 137
rect 183 136 184 137
rect 184 136 185 137
rect 185 136 186 137
rect 186 136 187 137
rect 187 136 188 137
rect 188 136 189 137
rect 189 136 190 137
rect 190 136 191 137
rect 191 136 192 137
rect 192 136 193 137
rect 193 136 194 137
rect 194 136 195 137
rect 195 136 196 137
rect 196 136 197 137
rect 197 136 198 137
rect 198 136 199 137
rect 199 136 200 137
rect 200 136 201 137
rect 201 136 202 137
rect 202 136 203 137
rect 203 136 204 137
rect 204 136 205 137
rect 205 136 206 137
rect 206 136 207 137
rect 207 136 208 137
rect 208 136 209 137
rect 209 136 210 137
rect 210 136 211 137
rect 211 136 212 137
rect 212 136 213 137
rect 213 136 214 137
rect 214 136 215 137
rect 215 136 216 137
rect 216 136 217 137
rect 217 136 218 137
rect 218 136 219 137
rect 219 136 220 137
rect 220 136 221 137
rect 240 136 241 137
rect 241 136 242 137
rect 242 136 243 137
rect 243 136 244 137
rect 244 136 245 137
rect 245 136 246 137
rect 246 136 247 137
rect 247 136 248 137
rect 248 136 249 137
rect 249 136 250 137
rect 250 136 251 137
rect 251 136 252 137
rect 252 136 253 137
rect 253 136 254 137
rect 254 136 255 137
rect 255 136 256 137
rect 256 136 257 137
rect 257 136 258 137
rect 258 136 259 137
rect 259 136 260 137
rect 260 136 261 137
rect 261 136 262 137
rect 262 136 263 137
rect 263 136 264 137
rect 264 136 265 137
rect 297 136 298 137
rect 298 136 299 137
rect 299 136 300 137
rect 300 136 301 137
rect 301 136 302 137
rect 307 136 308 137
rect 308 136 309 137
rect 309 136 310 137
rect 310 136 311 137
rect 311 136 312 137
rect 312 136 313 137
rect 313 136 314 137
rect 323 136 324 137
rect 324 136 325 137
rect 325 136 326 137
rect 326 136 327 137
rect 327 136 328 137
rect 328 136 329 137
rect 329 136 330 137
rect 330 136 331 137
rect 331 136 332 137
rect 332 136 333 137
rect 333 136 334 137
rect 334 136 335 137
rect 335 136 336 137
rect 336 136 337 137
rect 337 136 338 137
rect 338 136 339 137
rect 339 136 340 137
rect 340 136 341 137
rect 341 136 342 137
rect 342 136 343 137
rect 343 136 344 137
rect 344 136 345 137
rect 345 136 346 137
rect 346 136 347 137
rect 347 136 348 137
rect 348 136 349 137
rect 370 136 371 137
rect 371 136 372 137
rect 372 136 373 137
rect 373 136 374 137
rect 374 136 375 137
rect 375 136 376 137
rect 376 136 377 137
rect 377 136 378 137
rect 182 135 183 136
rect 183 135 184 136
rect 184 135 185 136
rect 185 135 186 136
rect 186 135 187 136
rect 187 135 188 136
rect 188 135 189 136
rect 189 135 190 136
rect 190 135 191 136
rect 191 135 192 136
rect 192 135 193 136
rect 193 135 194 136
rect 194 135 195 136
rect 195 135 196 136
rect 196 135 197 136
rect 197 135 198 136
rect 198 135 199 136
rect 199 135 200 136
rect 200 135 201 136
rect 201 135 202 136
rect 202 135 203 136
rect 203 135 204 136
rect 204 135 205 136
rect 205 135 206 136
rect 206 135 207 136
rect 207 135 208 136
rect 208 135 209 136
rect 209 135 210 136
rect 210 135 211 136
rect 211 135 212 136
rect 212 135 213 136
rect 213 135 214 136
rect 214 135 215 136
rect 215 135 216 136
rect 216 135 217 136
rect 217 135 218 136
rect 218 135 219 136
rect 219 135 220 136
rect 220 135 221 136
rect 221 135 222 136
rect 222 135 223 136
rect 223 135 224 136
rect 224 135 225 136
rect 225 135 226 136
rect 226 135 227 136
rect 227 135 228 136
rect 232 135 233 136
rect 233 135 234 136
rect 234 135 235 136
rect 235 135 236 136
rect 236 135 237 136
rect 237 135 238 136
rect 238 135 239 136
rect 239 135 240 136
rect 240 135 241 136
rect 241 135 242 136
rect 242 135 243 136
rect 243 135 244 136
rect 244 135 245 136
rect 245 135 246 136
rect 246 135 247 136
rect 247 135 248 136
rect 248 135 249 136
rect 249 135 250 136
rect 250 135 251 136
rect 251 135 252 136
rect 252 135 253 136
rect 253 135 254 136
rect 254 135 255 136
rect 255 135 256 136
rect 256 135 257 136
rect 257 135 258 136
rect 258 135 259 136
rect 259 135 260 136
rect 260 135 261 136
rect 261 135 262 136
rect 262 135 263 136
rect 296 135 297 136
rect 297 135 298 136
rect 298 135 299 136
rect 299 135 300 136
rect 300 135 301 136
rect 307 135 308 136
rect 308 135 309 136
rect 309 135 310 136
rect 310 135 311 136
rect 311 135 312 136
rect 312 135 313 136
rect 313 135 314 136
rect 326 135 327 136
rect 327 135 328 136
rect 328 135 329 136
rect 329 135 330 136
rect 330 135 331 136
rect 331 135 332 136
rect 332 135 333 136
rect 333 135 334 136
rect 334 135 335 136
rect 335 135 336 136
rect 336 135 337 136
rect 337 135 338 136
rect 338 135 339 136
rect 339 135 340 136
rect 340 135 341 136
rect 341 135 342 136
rect 342 135 343 136
rect 343 135 344 136
rect 344 135 345 136
rect 345 135 346 136
rect 346 135 347 136
rect 347 135 348 136
rect 348 135 349 136
rect 349 135 350 136
rect 350 135 351 136
rect 351 135 352 136
rect 352 135 353 136
rect 370 135 371 136
rect 371 135 372 136
rect 372 135 373 136
rect 373 135 374 136
rect 374 135 375 136
rect 375 135 376 136
rect 376 135 377 136
rect 377 135 378 136
rect 183 134 184 135
rect 184 134 185 135
rect 185 134 186 135
rect 186 134 187 135
rect 187 134 188 135
rect 188 134 189 135
rect 189 134 190 135
rect 190 134 191 135
rect 191 134 192 135
rect 192 134 193 135
rect 193 134 194 135
rect 194 134 195 135
rect 195 134 196 135
rect 196 134 197 135
rect 197 134 198 135
rect 198 134 199 135
rect 199 134 200 135
rect 200 134 201 135
rect 201 134 202 135
rect 202 134 203 135
rect 203 134 204 135
rect 204 134 205 135
rect 205 134 206 135
rect 206 134 207 135
rect 207 134 208 135
rect 208 134 209 135
rect 209 134 210 135
rect 210 134 211 135
rect 211 134 212 135
rect 212 134 213 135
rect 213 134 214 135
rect 214 134 215 135
rect 215 134 216 135
rect 216 134 217 135
rect 217 134 218 135
rect 218 134 219 135
rect 219 134 220 135
rect 220 134 221 135
rect 221 134 222 135
rect 222 134 223 135
rect 223 134 224 135
rect 224 134 225 135
rect 225 134 226 135
rect 226 134 227 135
rect 227 134 228 135
rect 228 134 229 135
rect 229 134 230 135
rect 230 134 231 135
rect 231 134 232 135
rect 232 134 233 135
rect 233 134 234 135
rect 234 134 235 135
rect 235 134 236 135
rect 236 134 237 135
rect 237 134 238 135
rect 238 134 239 135
rect 239 134 240 135
rect 240 134 241 135
rect 241 134 242 135
rect 242 134 243 135
rect 243 134 244 135
rect 244 134 245 135
rect 245 134 246 135
rect 246 134 247 135
rect 247 134 248 135
rect 248 134 249 135
rect 249 134 250 135
rect 250 134 251 135
rect 251 134 252 135
rect 252 134 253 135
rect 253 134 254 135
rect 254 134 255 135
rect 255 134 256 135
rect 256 134 257 135
rect 257 134 258 135
rect 258 134 259 135
rect 259 134 260 135
rect 260 134 261 135
rect 261 134 262 135
rect 295 134 296 135
rect 296 134 297 135
rect 297 134 298 135
rect 298 134 299 135
rect 299 134 300 135
rect 307 134 308 135
rect 308 134 309 135
rect 309 134 310 135
rect 310 134 311 135
rect 311 134 312 135
rect 312 134 313 135
rect 313 134 314 135
rect 329 134 330 135
rect 330 134 331 135
rect 331 134 332 135
rect 332 134 333 135
rect 333 134 334 135
rect 334 134 335 135
rect 335 134 336 135
rect 336 134 337 135
rect 337 134 338 135
rect 338 134 339 135
rect 339 134 340 135
rect 340 134 341 135
rect 341 134 342 135
rect 342 134 343 135
rect 343 134 344 135
rect 344 134 345 135
rect 345 134 346 135
rect 346 134 347 135
rect 347 134 348 135
rect 348 134 349 135
rect 349 134 350 135
rect 350 134 351 135
rect 351 134 352 135
rect 352 134 353 135
rect 353 134 354 135
rect 354 134 355 135
rect 355 134 356 135
rect 370 134 371 135
rect 371 134 372 135
rect 372 134 373 135
rect 373 134 374 135
rect 374 134 375 135
rect 375 134 376 135
rect 376 134 377 135
rect 377 134 378 135
rect 184 133 185 134
rect 185 133 186 134
rect 186 133 187 134
rect 187 133 188 134
rect 188 133 189 134
rect 189 133 190 134
rect 190 133 191 134
rect 191 133 192 134
rect 192 133 193 134
rect 193 133 194 134
rect 194 133 195 134
rect 195 133 196 134
rect 196 133 197 134
rect 197 133 198 134
rect 198 133 199 134
rect 199 133 200 134
rect 200 133 201 134
rect 201 133 202 134
rect 202 133 203 134
rect 203 133 204 134
rect 204 133 205 134
rect 205 133 206 134
rect 206 133 207 134
rect 207 133 208 134
rect 208 133 209 134
rect 209 133 210 134
rect 210 133 211 134
rect 211 133 212 134
rect 212 133 213 134
rect 213 133 214 134
rect 214 133 215 134
rect 215 133 216 134
rect 216 133 217 134
rect 217 133 218 134
rect 218 133 219 134
rect 219 133 220 134
rect 220 133 221 134
rect 221 133 222 134
rect 222 133 223 134
rect 223 133 224 134
rect 224 133 225 134
rect 225 133 226 134
rect 226 133 227 134
rect 227 133 228 134
rect 228 133 229 134
rect 229 133 230 134
rect 230 133 231 134
rect 231 133 232 134
rect 232 133 233 134
rect 233 133 234 134
rect 234 133 235 134
rect 235 133 236 134
rect 236 133 237 134
rect 237 133 238 134
rect 238 133 239 134
rect 239 133 240 134
rect 240 133 241 134
rect 241 133 242 134
rect 242 133 243 134
rect 243 133 244 134
rect 244 133 245 134
rect 245 133 246 134
rect 246 133 247 134
rect 247 133 248 134
rect 248 133 249 134
rect 249 133 250 134
rect 250 133 251 134
rect 251 133 252 134
rect 252 133 253 134
rect 253 133 254 134
rect 254 133 255 134
rect 255 133 256 134
rect 256 133 257 134
rect 257 133 258 134
rect 258 133 259 134
rect 259 133 260 134
rect 294 133 295 134
rect 295 133 296 134
rect 296 133 297 134
rect 297 133 298 134
rect 298 133 299 134
rect 299 133 300 134
rect 307 133 308 134
rect 308 133 309 134
rect 309 133 310 134
rect 310 133 311 134
rect 311 133 312 134
rect 312 133 313 134
rect 313 133 314 134
rect 332 133 333 134
rect 333 133 334 134
rect 334 133 335 134
rect 335 133 336 134
rect 336 133 337 134
rect 337 133 338 134
rect 338 133 339 134
rect 339 133 340 134
rect 340 133 341 134
rect 341 133 342 134
rect 342 133 343 134
rect 343 133 344 134
rect 344 133 345 134
rect 345 133 346 134
rect 346 133 347 134
rect 347 133 348 134
rect 348 133 349 134
rect 349 133 350 134
rect 350 133 351 134
rect 351 133 352 134
rect 352 133 353 134
rect 353 133 354 134
rect 354 133 355 134
rect 355 133 356 134
rect 356 133 357 134
rect 357 133 358 134
rect 358 133 359 134
rect 369 133 370 134
rect 370 133 371 134
rect 371 133 372 134
rect 372 133 373 134
rect 373 133 374 134
rect 374 133 375 134
rect 375 133 376 134
rect 376 133 377 134
rect 185 132 186 133
rect 186 132 187 133
rect 187 132 188 133
rect 188 132 189 133
rect 189 132 190 133
rect 190 132 191 133
rect 191 132 192 133
rect 192 132 193 133
rect 193 132 194 133
rect 194 132 195 133
rect 195 132 196 133
rect 196 132 197 133
rect 197 132 198 133
rect 198 132 199 133
rect 199 132 200 133
rect 200 132 201 133
rect 201 132 202 133
rect 202 132 203 133
rect 203 132 204 133
rect 204 132 205 133
rect 205 132 206 133
rect 206 132 207 133
rect 207 132 208 133
rect 208 132 209 133
rect 209 132 210 133
rect 210 132 211 133
rect 211 132 212 133
rect 212 132 213 133
rect 213 132 214 133
rect 214 132 215 133
rect 215 132 216 133
rect 216 132 217 133
rect 217 132 218 133
rect 218 132 219 133
rect 219 132 220 133
rect 220 132 221 133
rect 221 132 222 133
rect 222 132 223 133
rect 223 132 224 133
rect 224 132 225 133
rect 225 132 226 133
rect 226 132 227 133
rect 227 132 228 133
rect 228 132 229 133
rect 229 132 230 133
rect 230 132 231 133
rect 231 132 232 133
rect 232 132 233 133
rect 233 132 234 133
rect 234 132 235 133
rect 235 132 236 133
rect 236 132 237 133
rect 237 132 238 133
rect 238 132 239 133
rect 239 132 240 133
rect 240 132 241 133
rect 241 132 242 133
rect 242 132 243 133
rect 243 132 244 133
rect 244 132 245 133
rect 245 132 246 133
rect 246 132 247 133
rect 247 132 248 133
rect 248 132 249 133
rect 249 132 250 133
rect 250 132 251 133
rect 251 132 252 133
rect 252 132 253 133
rect 253 132 254 133
rect 254 132 255 133
rect 255 132 256 133
rect 256 132 257 133
rect 257 132 258 133
rect 294 132 295 133
rect 295 132 296 133
rect 296 132 297 133
rect 297 132 298 133
rect 298 132 299 133
rect 307 132 308 133
rect 308 132 309 133
rect 309 132 310 133
rect 310 132 311 133
rect 311 132 312 133
rect 312 132 313 133
rect 313 132 314 133
rect 336 132 337 133
rect 337 132 338 133
rect 338 132 339 133
rect 339 132 340 133
rect 340 132 341 133
rect 341 132 342 133
rect 342 132 343 133
rect 343 132 344 133
rect 344 132 345 133
rect 345 132 346 133
rect 346 132 347 133
rect 347 132 348 133
rect 348 132 349 133
rect 349 132 350 133
rect 350 132 351 133
rect 351 132 352 133
rect 352 132 353 133
rect 353 132 354 133
rect 354 132 355 133
rect 355 132 356 133
rect 356 132 357 133
rect 357 132 358 133
rect 358 132 359 133
rect 359 132 360 133
rect 360 132 361 133
rect 361 132 362 133
rect 362 132 363 133
rect 367 132 368 133
rect 368 132 369 133
rect 369 132 370 133
rect 370 132 371 133
rect 371 132 372 133
rect 372 132 373 133
rect 373 132 374 133
rect 374 132 375 133
rect 375 132 376 133
rect 376 132 377 133
rect 186 131 187 132
rect 187 131 188 132
rect 188 131 189 132
rect 189 131 190 132
rect 190 131 191 132
rect 191 131 192 132
rect 192 131 193 132
rect 193 131 194 132
rect 195 131 196 132
rect 196 131 197 132
rect 197 131 198 132
rect 198 131 199 132
rect 199 131 200 132
rect 200 131 201 132
rect 201 131 202 132
rect 202 131 203 132
rect 203 131 204 132
rect 204 131 205 132
rect 205 131 206 132
rect 206 131 207 132
rect 207 131 208 132
rect 208 131 209 132
rect 209 131 210 132
rect 210 131 211 132
rect 211 131 212 132
rect 212 131 213 132
rect 213 131 214 132
rect 214 131 215 132
rect 215 131 216 132
rect 216 131 217 132
rect 217 131 218 132
rect 218 131 219 132
rect 219 131 220 132
rect 220 131 221 132
rect 221 131 222 132
rect 222 131 223 132
rect 223 131 224 132
rect 224 131 225 132
rect 225 131 226 132
rect 226 131 227 132
rect 227 131 228 132
rect 228 131 229 132
rect 229 131 230 132
rect 230 131 231 132
rect 231 131 232 132
rect 232 131 233 132
rect 233 131 234 132
rect 234 131 235 132
rect 235 131 236 132
rect 236 131 237 132
rect 237 131 238 132
rect 238 131 239 132
rect 239 131 240 132
rect 240 131 241 132
rect 241 131 242 132
rect 242 131 243 132
rect 243 131 244 132
rect 244 131 245 132
rect 245 131 246 132
rect 246 131 247 132
rect 247 131 248 132
rect 248 131 249 132
rect 249 131 250 132
rect 250 131 251 132
rect 251 131 252 132
rect 252 131 253 132
rect 253 131 254 132
rect 254 131 255 132
rect 255 131 256 132
rect 256 131 257 132
rect 293 131 294 132
rect 294 131 295 132
rect 295 131 296 132
rect 296 131 297 132
rect 297 131 298 132
rect 307 131 308 132
rect 308 131 309 132
rect 309 131 310 132
rect 310 131 311 132
rect 311 131 312 132
rect 312 131 313 132
rect 313 131 314 132
rect 340 131 341 132
rect 341 131 342 132
rect 342 131 343 132
rect 343 131 344 132
rect 344 131 345 132
rect 345 131 346 132
rect 346 131 347 132
rect 347 131 348 132
rect 348 131 349 132
rect 349 131 350 132
rect 350 131 351 132
rect 351 131 352 132
rect 352 131 353 132
rect 353 131 354 132
rect 354 131 355 132
rect 355 131 356 132
rect 356 131 357 132
rect 357 131 358 132
rect 358 131 359 132
rect 359 131 360 132
rect 360 131 361 132
rect 361 131 362 132
rect 362 131 363 132
rect 363 131 364 132
rect 364 131 365 132
rect 365 131 366 132
rect 366 131 367 132
rect 367 131 368 132
rect 368 131 369 132
rect 369 131 370 132
rect 370 131 371 132
rect 371 131 372 132
rect 372 131 373 132
rect 373 131 374 132
rect 374 131 375 132
rect 375 131 376 132
rect 186 130 187 131
rect 187 130 188 131
rect 188 130 189 131
rect 189 130 190 131
rect 190 130 191 131
rect 191 130 192 131
rect 192 130 193 131
rect 193 130 194 131
rect 199 130 200 131
rect 200 130 201 131
rect 201 130 202 131
rect 202 130 203 131
rect 203 130 204 131
rect 204 130 205 131
rect 205 130 206 131
rect 206 130 207 131
rect 207 130 208 131
rect 208 130 209 131
rect 209 130 210 131
rect 210 130 211 131
rect 211 130 212 131
rect 212 130 213 131
rect 213 130 214 131
rect 214 130 215 131
rect 215 130 216 131
rect 216 130 217 131
rect 217 130 218 131
rect 218 130 219 131
rect 219 130 220 131
rect 220 130 221 131
rect 221 130 222 131
rect 222 130 223 131
rect 223 130 224 131
rect 224 130 225 131
rect 225 130 226 131
rect 226 130 227 131
rect 227 130 228 131
rect 228 130 229 131
rect 229 130 230 131
rect 230 130 231 131
rect 231 130 232 131
rect 232 130 233 131
rect 233 130 234 131
rect 234 130 235 131
rect 235 130 236 131
rect 236 130 237 131
rect 237 130 238 131
rect 238 130 239 131
rect 239 130 240 131
rect 240 130 241 131
rect 241 130 242 131
rect 242 130 243 131
rect 243 130 244 131
rect 244 130 245 131
rect 245 130 246 131
rect 246 130 247 131
rect 247 130 248 131
rect 248 130 249 131
rect 249 130 250 131
rect 250 130 251 131
rect 251 130 252 131
rect 252 130 253 131
rect 253 130 254 131
rect 254 130 255 131
rect 292 130 293 131
rect 293 130 294 131
rect 294 130 295 131
rect 295 130 296 131
rect 296 130 297 131
rect 306 130 307 131
rect 307 130 308 131
rect 308 130 309 131
rect 309 130 310 131
rect 310 130 311 131
rect 311 130 312 131
rect 312 130 313 131
rect 344 130 345 131
rect 345 130 346 131
rect 346 130 347 131
rect 347 130 348 131
rect 348 130 349 131
rect 349 130 350 131
rect 350 130 351 131
rect 351 130 352 131
rect 352 130 353 131
rect 353 130 354 131
rect 354 130 355 131
rect 355 130 356 131
rect 356 130 357 131
rect 357 130 358 131
rect 358 130 359 131
rect 359 130 360 131
rect 360 130 361 131
rect 361 130 362 131
rect 362 130 363 131
rect 363 130 364 131
rect 364 130 365 131
rect 365 130 366 131
rect 366 130 367 131
rect 367 130 368 131
rect 368 130 369 131
rect 369 130 370 131
rect 370 130 371 131
rect 371 130 372 131
rect 372 130 373 131
rect 373 130 374 131
rect 374 130 375 131
rect 375 130 376 131
rect 186 129 187 130
rect 187 129 188 130
rect 188 129 189 130
rect 189 129 190 130
rect 190 129 191 130
rect 191 129 192 130
rect 192 129 193 130
rect 193 129 194 130
rect 203 129 204 130
rect 204 129 205 130
rect 205 129 206 130
rect 206 129 207 130
rect 207 129 208 130
rect 208 129 209 130
rect 209 129 210 130
rect 210 129 211 130
rect 211 129 212 130
rect 212 129 213 130
rect 213 129 214 130
rect 214 129 215 130
rect 215 129 216 130
rect 216 129 217 130
rect 217 129 218 130
rect 218 129 219 130
rect 219 129 220 130
rect 220 129 221 130
rect 221 129 222 130
rect 222 129 223 130
rect 223 129 224 130
rect 224 129 225 130
rect 225 129 226 130
rect 226 129 227 130
rect 227 129 228 130
rect 228 129 229 130
rect 229 129 230 130
rect 230 129 231 130
rect 231 129 232 130
rect 232 129 233 130
rect 233 129 234 130
rect 234 129 235 130
rect 235 129 236 130
rect 236 129 237 130
rect 237 129 238 130
rect 238 129 239 130
rect 239 129 240 130
rect 240 129 241 130
rect 241 129 242 130
rect 242 129 243 130
rect 243 129 244 130
rect 244 129 245 130
rect 245 129 246 130
rect 246 129 247 130
rect 247 129 248 130
rect 248 129 249 130
rect 249 129 250 130
rect 250 129 251 130
rect 251 129 252 130
rect 291 129 292 130
rect 292 129 293 130
rect 293 129 294 130
rect 294 129 295 130
rect 295 129 296 130
rect 296 129 297 130
rect 306 129 307 130
rect 307 129 308 130
rect 308 129 309 130
rect 309 129 310 130
rect 310 129 311 130
rect 311 129 312 130
rect 312 129 313 130
rect 348 129 349 130
rect 349 129 350 130
rect 350 129 351 130
rect 351 129 352 130
rect 352 129 353 130
rect 353 129 354 130
rect 354 129 355 130
rect 355 129 356 130
rect 356 129 357 130
rect 357 129 358 130
rect 358 129 359 130
rect 359 129 360 130
rect 360 129 361 130
rect 361 129 362 130
rect 362 129 363 130
rect 363 129 364 130
rect 364 129 365 130
rect 365 129 366 130
rect 366 129 367 130
rect 367 129 368 130
rect 368 129 369 130
rect 369 129 370 130
rect 370 129 371 130
rect 371 129 372 130
rect 372 129 373 130
rect 373 129 374 130
rect 374 129 375 130
rect 186 128 187 129
rect 187 128 188 129
rect 188 128 189 129
rect 189 128 190 129
rect 190 128 191 129
rect 191 128 192 129
rect 192 128 193 129
rect 193 128 194 129
rect 207 128 208 129
rect 208 128 209 129
rect 209 128 210 129
rect 210 128 211 129
rect 211 128 212 129
rect 212 128 213 129
rect 213 128 214 129
rect 214 128 215 129
rect 215 128 216 129
rect 216 128 217 129
rect 217 128 218 129
rect 218 128 219 129
rect 219 128 220 129
rect 220 128 221 129
rect 221 128 222 129
rect 222 128 223 129
rect 223 128 224 129
rect 224 128 225 129
rect 225 128 226 129
rect 226 128 227 129
rect 227 128 228 129
rect 228 128 229 129
rect 229 128 230 129
rect 230 128 231 129
rect 231 128 232 129
rect 232 128 233 129
rect 233 128 234 129
rect 234 128 235 129
rect 235 128 236 129
rect 236 128 237 129
rect 237 128 238 129
rect 238 128 239 129
rect 239 128 240 129
rect 240 128 241 129
rect 241 128 242 129
rect 242 128 243 129
rect 243 128 244 129
rect 244 128 245 129
rect 245 128 246 129
rect 246 128 247 129
rect 247 128 248 129
rect 248 128 249 129
rect 249 128 250 129
rect 291 128 292 129
rect 292 128 293 129
rect 293 128 294 129
rect 294 128 295 129
rect 295 128 296 129
rect 306 128 307 129
rect 307 128 308 129
rect 308 128 309 129
rect 309 128 310 129
rect 310 128 311 129
rect 311 128 312 129
rect 312 128 313 129
rect 351 128 352 129
rect 352 128 353 129
rect 353 128 354 129
rect 354 128 355 129
rect 355 128 356 129
rect 356 128 357 129
rect 357 128 358 129
rect 358 128 359 129
rect 359 128 360 129
rect 360 128 361 129
rect 361 128 362 129
rect 362 128 363 129
rect 363 128 364 129
rect 364 128 365 129
rect 365 128 366 129
rect 366 128 367 129
rect 367 128 368 129
rect 368 128 369 129
rect 369 128 370 129
rect 370 128 371 129
rect 371 128 372 129
rect 372 128 373 129
rect 373 128 374 129
rect 187 127 188 128
rect 188 127 189 128
rect 189 127 190 128
rect 190 127 191 128
rect 191 127 192 128
rect 192 127 193 128
rect 193 127 194 128
rect 212 127 213 128
rect 213 127 214 128
rect 214 127 215 128
rect 215 127 216 128
rect 216 127 217 128
rect 217 127 218 128
rect 218 127 219 128
rect 219 127 220 128
rect 220 127 221 128
rect 221 127 222 128
rect 222 127 223 128
rect 223 127 224 128
rect 224 127 225 128
rect 225 127 226 128
rect 226 127 227 128
rect 227 127 228 128
rect 228 127 229 128
rect 229 127 230 128
rect 230 127 231 128
rect 231 127 232 128
rect 232 127 233 128
rect 233 127 234 128
rect 234 127 235 128
rect 235 127 236 128
rect 236 127 237 128
rect 237 127 238 128
rect 238 127 239 128
rect 239 127 240 128
rect 240 127 241 128
rect 241 127 242 128
rect 242 127 243 128
rect 243 127 244 128
rect 244 127 245 128
rect 245 127 246 128
rect 246 127 247 128
rect 290 127 291 128
rect 291 127 292 128
rect 292 127 293 128
rect 293 127 294 128
rect 294 127 295 128
rect 306 127 307 128
rect 307 127 308 128
rect 308 127 309 128
rect 309 127 310 128
rect 310 127 311 128
rect 311 127 312 128
rect 312 127 313 128
rect 354 127 355 128
rect 355 127 356 128
rect 356 127 357 128
rect 357 127 358 128
rect 358 127 359 128
rect 359 127 360 128
rect 360 127 361 128
rect 361 127 362 128
rect 362 127 363 128
rect 363 127 364 128
rect 364 127 365 128
rect 365 127 366 128
rect 366 127 367 128
rect 367 127 368 128
rect 368 127 369 128
rect 369 127 370 128
rect 370 127 371 128
rect 371 127 372 128
rect 187 126 188 127
rect 188 126 189 127
rect 189 126 190 127
rect 190 126 191 127
rect 191 126 192 127
rect 192 126 193 127
rect 193 126 194 127
rect 218 126 219 127
rect 219 126 220 127
rect 220 126 221 127
rect 221 126 222 127
rect 222 126 223 127
rect 223 126 224 127
rect 224 126 225 127
rect 225 126 226 127
rect 226 126 227 127
rect 227 126 228 127
rect 228 126 229 127
rect 229 126 230 127
rect 230 126 231 127
rect 231 126 232 127
rect 232 126 233 127
rect 233 126 234 127
rect 234 126 235 127
rect 235 126 236 127
rect 236 126 237 127
rect 237 126 238 127
rect 238 126 239 127
rect 239 126 240 127
rect 240 126 241 127
rect 241 126 242 127
rect 289 126 290 127
rect 290 126 291 127
rect 291 126 292 127
rect 292 126 293 127
rect 293 126 294 127
rect 305 126 306 127
rect 306 126 307 127
rect 307 126 308 127
rect 308 126 309 127
rect 309 126 310 127
rect 310 126 311 127
rect 311 126 312 127
rect 312 126 313 127
rect 358 126 359 127
rect 359 126 360 127
rect 360 126 361 127
rect 361 126 362 127
rect 362 126 363 127
rect 363 126 364 127
rect 364 126 365 127
rect 365 126 366 127
rect 366 126 367 127
rect 367 126 368 127
rect 368 126 369 127
rect 369 126 370 127
rect 187 125 188 126
rect 188 125 189 126
rect 189 125 190 126
rect 190 125 191 126
rect 191 125 192 126
rect 192 125 193 126
rect 193 125 194 126
rect 194 125 195 126
rect 288 125 289 126
rect 289 125 290 126
rect 290 125 291 126
rect 291 125 292 126
rect 292 125 293 126
rect 305 125 306 126
rect 306 125 307 126
rect 307 125 308 126
rect 308 125 309 126
rect 309 125 310 126
rect 310 125 311 126
rect 311 125 312 126
rect 312 125 313 126
rect 363 125 364 126
rect 364 125 365 126
rect 365 125 366 126
rect 187 124 188 125
rect 188 124 189 125
rect 189 124 190 125
rect 190 124 191 125
rect 191 124 192 125
rect 192 124 193 125
rect 193 124 194 125
rect 194 124 195 125
rect 287 124 288 125
rect 288 124 289 125
rect 289 124 290 125
rect 290 124 291 125
rect 291 124 292 125
rect 305 124 306 125
rect 306 124 307 125
rect 307 124 308 125
rect 308 124 309 125
rect 309 124 310 125
rect 310 124 311 125
rect 311 124 312 125
rect 187 123 188 124
rect 188 123 189 124
rect 189 123 190 124
rect 190 123 191 124
rect 191 123 192 124
rect 192 123 193 124
rect 193 123 194 124
rect 194 123 195 124
rect 287 123 288 124
rect 288 123 289 124
rect 289 123 290 124
rect 290 123 291 124
rect 304 123 305 124
rect 305 123 306 124
rect 306 123 307 124
rect 307 123 308 124
rect 308 123 309 124
rect 309 123 310 124
rect 310 123 311 124
rect 311 123 312 124
rect 188 122 189 123
rect 189 122 190 123
rect 190 122 191 123
rect 191 122 192 123
rect 192 122 193 123
rect 193 122 194 123
rect 194 122 195 123
rect 286 122 287 123
rect 287 122 288 123
rect 288 122 289 123
rect 289 122 290 123
rect 290 122 291 123
rect 304 122 305 123
rect 305 122 306 123
rect 306 122 307 123
rect 307 122 308 123
rect 308 122 309 123
rect 309 122 310 123
rect 310 122 311 123
rect 311 122 312 123
rect 188 121 189 122
rect 189 121 190 122
rect 190 121 191 122
rect 191 121 192 122
rect 192 121 193 122
rect 193 121 194 122
rect 194 121 195 122
rect 285 121 286 122
rect 286 121 287 122
rect 287 121 288 122
rect 288 121 289 122
rect 289 121 290 122
rect 303 121 304 122
rect 304 121 305 122
rect 305 121 306 122
rect 306 121 307 122
rect 307 121 308 122
rect 308 121 309 122
rect 309 121 310 122
rect 310 121 311 122
rect 326 121 327 122
rect 327 121 328 122
rect 328 121 329 122
rect 329 121 330 122
rect 330 121 331 122
rect 188 120 189 121
rect 189 120 190 121
rect 190 120 191 121
rect 191 120 192 121
rect 192 120 193 121
rect 193 120 194 121
rect 194 120 195 121
rect 195 120 196 121
rect 284 120 285 121
rect 285 120 286 121
rect 286 120 287 121
rect 287 120 288 121
rect 303 120 304 121
rect 304 120 305 121
rect 305 120 306 121
rect 306 120 307 121
rect 307 120 308 121
rect 308 120 309 121
rect 309 120 310 121
rect 310 120 311 121
rect 324 120 325 121
rect 325 120 326 121
rect 326 120 327 121
rect 327 120 328 121
rect 328 120 329 121
rect 329 120 330 121
rect 330 120 331 121
rect 331 120 332 121
rect 332 120 333 121
rect 189 119 190 120
rect 190 119 191 120
rect 191 119 192 120
rect 192 119 193 120
rect 193 119 194 120
rect 194 119 195 120
rect 195 119 196 120
rect 283 119 284 120
rect 284 119 285 120
rect 285 119 286 120
rect 286 119 287 120
rect 302 119 303 120
rect 303 119 304 120
rect 304 119 305 120
rect 305 119 306 120
rect 306 119 307 120
rect 307 119 308 120
rect 308 119 309 120
rect 309 119 310 120
rect 310 119 311 120
rect 323 119 324 120
rect 324 119 325 120
rect 325 119 326 120
rect 332 119 333 120
rect 333 119 334 120
rect 334 119 335 120
rect 189 118 190 119
rect 190 118 191 119
rect 191 118 192 119
rect 192 118 193 119
rect 193 118 194 119
rect 194 118 195 119
rect 195 118 196 119
rect 283 118 284 119
rect 284 118 285 119
rect 285 118 286 119
rect 301 118 302 119
rect 302 118 303 119
rect 303 118 304 119
rect 304 118 305 119
rect 305 118 306 119
rect 306 118 307 119
rect 307 118 308 119
rect 308 118 309 119
rect 309 118 310 119
rect 322 118 323 119
rect 323 118 324 119
rect 333 118 334 119
rect 334 118 335 119
rect 335 118 336 119
rect 189 117 190 118
rect 190 117 191 118
rect 191 117 192 118
rect 192 117 193 118
rect 193 117 194 118
rect 194 117 195 118
rect 195 117 196 118
rect 282 117 283 118
rect 283 117 284 118
rect 284 117 285 118
rect 300 117 301 118
rect 301 117 302 118
rect 302 117 303 118
rect 303 117 304 118
rect 304 117 305 118
rect 305 117 306 118
rect 306 117 307 118
rect 307 117 308 118
rect 308 117 309 118
rect 321 117 322 118
rect 322 117 323 118
rect 323 117 324 118
rect 325 117 326 118
rect 326 117 327 118
rect 327 117 328 118
rect 328 117 329 118
rect 329 117 330 118
rect 330 117 331 118
rect 331 117 332 118
rect 334 117 335 118
rect 335 117 336 118
rect 189 116 190 117
rect 190 116 191 117
rect 191 116 192 117
rect 192 116 193 117
rect 193 116 194 117
rect 194 116 195 117
rect 195 116 196 117
rect 196 116 197 117
rect 281 116 282 117
rect 282 116 283 117
rect 283 116 284 117
rect 300 116 301 117
rect 301 116 302 117
rect 302 116 303 117
rect 303 116 304 117
rect 304 116 305 117
rect 305 116 306 117
rect 306 116 307 117
rect 307 116 308 117
rect 308 116 309 117
rect 321 116 322 117
rect 322 116 323 117
rect 325 116 326 117
rect 326 116 327 117
rect 327 116 328 117
rect 328 116 329 117
rect 329 116 330 117
rect 330 116 331 117
rect 331 116 332 117
rect 335 116 336 117
rect 336 116 337 117
rect 190 115 191 116
rect 191 115 192 116
rect 192 115 193 116
rect 193 115 194 116
rect 194 115 195 116
rect 195 115 196 116
rect 196 115 197 116
rect 281 115 282 116
rect 299 115 300 116
rect 300 115 301 116
rect 301 115 302 116
rect 302 115 303 116
rect 303 115 304 116
rect 304 115 305 116
rect 305 115 306 116
rect 306 115 307 116
rect 307 115 308 116
rect 321 115 322 116
rect 322 115 323 116
rect 325 115 326 116
rect 326 115 327 116
rect 327 115 328 116
rect 331 115 332 116
rect 332 115 333 116
rect 335 115 336 116
rect 336 115 337 116
rect 190 114 191 115
rect 191 114 192 115
rect 192 114 193 115
rect 193 114 194 115
rect 194 114 195 115
rect 195 114 196 115
rect 196 114 197 115
rect 298 114 299 115
rect 299 114 300 115
rect 300 114 301 115
rect 301 114 302 115
rect 302 114 303 115
rect 303 114 304 115
rect 304 114 305 115
rect 305 114 306 115
rect 306 114 307 115
rect 321 114 322 115
rect 325 114 326 115
rect 326 114 327 115
rect 327 114 328 115
rect 330 114 331 115
rect 331 114 332 115
rect 335 114 336 115
rect 336 114 337 115
rect 190 113 191 114
rect 191 113 192 114
rect 192 113 193 114
rect 193 113 194 114
rect 194 113 195 114
rect 195 113 196 114
rect 196 113 197 114
rect 298 113 299 114
rect 299 113 300 114
rect 300 113 301 114
rect 301 113 302 114
rect 302 113 303 114
rect 303 113 304 114
rect 304 113 305 114
rect 305 113 306 114
rect 306 113 307 114
rect 320 113 321 114
rect 321 113 322 114
rect 325 113 326 114
rect 326 113 327 114
rect 327 113 328 114
rect 328 113 329 114
rect 329 113 330 114
rect 330 113 331 114
rect 331 113 332 114
rect 335 113 336 114
rect 336 113 337 114
rect 190 112 191 113
rect 191 112 192 113
rect 192 112 193 113
rect 193 112 194 113
rect 194 112 195 113
rect 195 112 196 113
rect 196 112 197 113
rect 197 112 198 113
rect 297 112 298 113
rect 298 112 299 113
rect 299 112 300 113
rect 300 112 301 113
rect 301 112 302 113
rect 302 112 303 113
rect 303 112 304 113
rect 304 112 305 113
rect 305 112 306 113
rect 321 112 322 113
rect 326 112 327 113
rect 327 112 328 113
rect 330 112 331 113
rect 331 112 332 113
rect 335 112 336 113
rect 336 112 337 113
rect 191 111 192 112
rect 192 111 193 112
rect 193 111 194 112
rect 194 111 195 112
rect 195 111 196 112
rect 196 111 197 112
rect 197 111 198 112
rect 296 111 297 112
rect 297 111 298 112
rect 298 111 299 112
rect 299 111 300 112
rect 300 111 301 112
rect 301 111 302 112
rect 302 111 303 112
rect 303 111 304 112
rect 304 111 305 112
rect 321 111 322 112
rect 322 111 323 112
rect 326 111 327 112
rect 327 111 328 112
rect 330 111 331 112
rect 331 111 332 112
rect 335 111 336 112
rect 336 111 337 112
rect 191 110 192 111
rect 192 110 193 111
rect 193 110 194 111
rect 194 110 195 111
rect 195 110 196 111
rect 196 110 197 111
rect 197 110 198 111
rect 295 110 296 111
rect 296 110 297 111
rect 297 110 298 111
rect 298 110 299 111
rect 299 110 300 111
rect 300 110 301 111
rect 301 110 302 111
rect 302 110 303 111
rect 303 110 304 111
rect 304 110 305 111
rect 321 110 322 111
rect 322 110 323 111
rect 326 110 327 111
rect 327 110 328 111
rect 330 110 331 111
rect 331 110 332 111
rect 332 110 333 111
rect 335 110 336 111
rect 336 110 337 111
rect 191 109 192 110
rect 192 109 193 110
rect 193 109 194 110
rect 194 109 195 110
rect 195 109 196 110
rect 196 109 197 110
rect 197 109 198 110
rect 198 109 199 110
rect 295 109 296 110
rect 296 109 297 110
rect 297 109 298 110
rect 298 109 299 110
rect 299 109 300 110
rect 300 109 301 110
rect 301 109 302 110
rect 302 109 303 110
rect 303 109 304 110
rect 322 109 323 110
rect 323 109 324 110
rect 326 109 327 110
rect 331 109 332 110
rect 334 109 335 110
rect 335 109 336 110
rect 192 108 193 109
rect 193 108 194 109
rect 194 108 195 109
rect 195 108 196 109
rect 196 108 197 109
rect 197 108 198 109
rect 198 108 199 109
rect 294 108 295 109
rect 295 108 296 109
rect 296 108 297 109
rect 297 108 298 109
rect 298 108 299 109
rect 299 108 300 109
rect 300 108 301 109
rect 301 108 302 109
rect 302 108 303 109
rect 322 108 323 109
rect 323 108 324 109
rect 324 108 325 109
rect 333 108 334 109
rect 334 108 335 109
rect 192 107 193 108
rect 193 107 194 108
rect 194 107 195 108
rect 195 107 196 108
rect 196 107 197 108
rect 197 107 198 108
rect 198 107 199 108
rect 293 107 294 108
rect 294 107 295 108
rect 295 107 296 108
rect 296 107 297 108
rect 297 107 298 108
rect 298 107 299 108
rect 299 107 300 108
rect 300 107 301 108
rect 301 107 302 108
rect 323 107 324 108
rect 324 107 325 108
rect 325 107 326 108
rect 331 107 332 108
rect 332 107 333 108
rect 333 107 334 108
rect 192 106 193 107
rect 193 106 194 107
rect 194 106 195 107
rect 195 106 196 107
rect 196 106 197 107
rect 197 106 198 107
rect 198 106 199 107
rect 199 106 200 107
rect 292 106 293 107
rect 293 106 294 107
rect 294 106 295 107
rect 295 106 296 107
rect 296 106 297 107
rect 297 106 298 107
rect 298 106 299 107
rect 299 106 300 107
rect 300 106 301 107
rect 301 106 302 107
rect 324 106 325 107
rect 325 106 326 107
rect 326 106 327 107
rect 327 106 328 107
rect 328 106 329 107
rect 329 106 330 107
rect 330 106 331 107
rect 331 106 332 107
rect 332 106 333 107
rect 192 105 193 106
rect 193 105 194 106
rect 194 105 195 106
rect 195 105 196 106
rect 196 105 197 106
rect 197 105 198 106
rect 198 105 199 106
rect 199 105 200 106
rect 292 105 293 106
rect 293 105 294 106
rect 294 105 295 106
rect 295 105 296 106
rect 296 105 297 106
rect 297 105 298 106
rect 298 105 299 106
rect 299 105 300 106
rect 300 105 301 106
rect 327 105 328 106
rect 328 105 329 106
rect 329 105 330 106
rect 330 105 331 106
rect 193 104 194 105
rect 194 104 195 105
rect 195 104 196 105
rect 196 104 197 105
rect 197 104 198 105
rect 198 104 199 105
rect 199 104 200 105
rect 291 104 292 105
rect 292 104 293 105
rect 293 104 294 105
rect 294 104 295 105
rect 295 104 296 105
rect 296 104 297 105
rect 297 104 298 105
rect 298 104 299 105
rect 299 104 300 105
rect 193 103 194 104
rect 194 103 195 104
rect 195 103 196 104
rect 196 103 197 104
rect 197 103 198 104
rect 198 103 199 104
rect 199 103 200 104
rect 200 103 201 104
rect 290 103 291 104
rect 291 103 292 104
rect 292 103 293 104
rect 293 103 294 104
rect 294 103 295 104
rect 295 103 296 104
rect 296 103 297 104
rect 297 103 298 104
rect 298 103 299 104
rect 193 102 194 103
rect 194 102 195 103
rect 195 102 196 103
rect 196 102 197 103
rect 197 102 198 103
rect 198 102 199 103
rect 199 102 200 103
rect 200 102 201 103
rect 289 102 290 103
rect 290 102 291 103
rect 291 102 292 103
rect 292 102 293 103
rect 293 102 294 103
rect 294 102 295 103
rect 295 102 296 103
rect 296 102 297 103
rect 297 102 298 103
rect 298 102 299 103
rect 194 101 195 102
rect 195 101 196 102
rect 196 101 197 102
rect 197 101 198 102
rect 198 101 199 102
rect 199 101 200 102
rect 200 101 201 102
rect 289 101 290 102
rect 290 101 291 102
rect 291 101 292 102
rect 292 101 293 102
rect 293 101 294 102
rect 294 101 295 102
rect 295 101 296 102
rect 296 101 297 102
rect 297 101 298 102
rect 194 100 195 101
rect 195 100 196 101
rect 196 100 197 101
rect 197 100 198 101
rect 198 100 199 101
rect 199 100 200 101
rect 200 100 201 101
rect 201 100 202 101
rect 288 100 289 101
rect 289 100 290 101
rect 290 100 291 101
rect 291 100 292 101
rect 292 100 293 101
rect 293 100 294 101
rect 294 100 295 101
rect 295 100 296 101
rect 296 100 297 101
rect 194 99 195 100
rect 195 99 196 100
rect 196 99 197 100
rect 197 99 198 100
rect 198 99 199 100
rect 199 99 200 100
rect 200 99 201 100
rect 201 99 202 100
rect 287 99 288 100
rect 288 99 289 100
rect 289 99 290 100
rect 290 99 291 100
rect 291 99 292 100
rect 292 99 293 100
rect 293 99 294 100
rect 294 99 295 100
rect 295 99 296 100
rect 296 99 297 100
rect 195 98 196 99
rect 196 98 197 99
rect 197 98 198 99
rect 198 98 199 99
rect 199 98 200 99
rect 200 98 201 99
rect 201 98 202 99
rect 202 98 203 99
rect 286 98 287 99
rect 287 98 288 99
rect 288 98 289 99
rect 289 98 290 99
rect 290 98 291 99
rect 291 98 292 99
rect 292 98 293 99
rect 293 98 294 99
rect 294 98 295 99
rect 295 98 296 99
rect 195 97 196 98
rect 196 97 197 98
rect 197 97 198 98
rect 198 97 199 98
rect 199 97 200 98
rect 200 97 201 98
rect 201 97 202 98
rect 202 97 203 98
rect 285 97 286 98
rect 286 97 287 98
rect 287 97 288 98
rect 288 97 289 98
rect 289 97 290 98
rect 290 97 291 98
rect 291 97 292 98
rect 292 97 293 98
rect 293 97 294 98
rect 294 97 295 98
rect 195 96 196 97
rect 196 96 197 97
rect 197 96 198 97
rect 198 96 199 97
rect 199 96 200 97
rect 200 96 201 97
rect 201 96 202 97
rect 202 96 203 97
rect 203 96 204 97
rect 285 96 286 97
rect 286 96 287 97
rect 287 96 288 97
rect 288 96 289 97
rect 289 96 290 97
rect 290 96 291 97
rect 291 96 292 97
rect 292 96 293 97
rect 293 96 294 97
rect 196 95 197 96
rect 197 95 198 96
rect 198 95 199 96
rect 199 95 200 96
rect 200 95 201 96
rect 201 95 202 96
rect 202 95 203 96
rect 203 95 204 96
rect 284 95 285 96
rect 285 95 286 96
rect 286 95 287 96
rect 287 95 288 96
rect 288 95 289 96
rect 289 95 290 96
rect 290 95 291 96
rect 291 95 292 96
rect 292 95 293 96
rect 196 94 197 95
rect 197 94 198 95
rect 198 94 199 95
rect 199 94 200 95
rect 200 94 201 95
rect 201 94 202 95
rect 202 94 203 95
rect 203 94 204 95
rect 204 94 205 95
rect 283 94 284 95
rect 284 94 285 95
rect 285 94 286 95
rect 286 94 287 95
rect 287 94 288 95
rect 288 94 289 95
rect 289 94 290 95
rect 290 94 291 95
rect 291 94 292 95
rect 292 94 293 95
rect 196 93 197 94
rect 197 93 198 94
rect 198 93 199 94
rect 199 93 200 94
rect 200 93 201 94
rect 201 93 202 94
rect 202 93 203 94
rect 203 93 204 94
rect 204 93 205 94
rect 282 93 283 94
rect 283 93 284 94
rect 284 93 285 94
rect 285 93 286 94
rect 286 93 287 94
rect 287 93 288 94
rect 288 93 289 94
rect 289 93 290 94
rect 290 93 291 94
rect 291 93 292 94
rect 197 92 198 93
rect 198 92 199 93
rect 199 92 200 93
rect 200 92 201 93
rect 201 92 202 93
rect 202 92 203 93
rect 203 92 204 93
rect 204 92 205 93
rect 205 92 206 93
rect 281 92 282 93
rect 282 92 283 93
rect 283 92 284 93
rect 284 92 285 93
rect 285 92 286 93
rect 286 92 287 93
rect 287 92 288 93
rect 288 92 289 93
rect 289 92 290 93
rect 290 92 291 93
rect 197 91 198 92
rect 198 91 199 92
rect 199 91 200 92
rect 200 91 201 92
rect 201 91 202 92
rect 202 91 203 92
rect 203 91 204 92
rect 204 91 205 92
rect 205 91 206 92
rect 206 91 207 92
rect 281 91 282 92
rect 282 91 283 92
rect 283 91 284 92
rect 284 91 285 92
rect 285 91 286 92
rect 286 91 287 92
rect 287 91 288 92
rect 288 91 289 92
rect 289 91 290 92
rect 198 90 199 91
rect 199 90 200 91
rect 200 90 201 91
rect 201 90 202 91
rect 202 90 203 91
rect 203 90 204 91
rect 204 90 205 91
rect 205 90 206 91
rect 206 90 207 91
rect 207 90 208 91
rect 280 90 281 91
rect 281 90 282 91
rect 282 90 283 91
rect 283 90 284 91
rect 284 90 285 91
rect 285 90 286 91
rect 286 90 287 91
rect 287 90 288 91
rect 288 90 289 91
rect 198 89 199 90
rect 199 89 200 90
rect 200 89 201 90
rect 201 89 202 90
rect 202 89 203 90
rect 203 89 204 90
rect 204 89 205 90
rect 205 89 206 90
rect 206 89 207 90
rect 207 89 208 90
rect 279 89 280 90
rect 280 89 281 90
rect 281 89 282 90
rect 282 89 283 90
rect 283 89 284 90
rect 284 89 285 90
rect 285 89 286 90
rect 286 89 287 90
rect 287 89 288 90
rect 288 89 289 90
rect 199 88 200 89
rect 200 88 201 89
rect 201 88 202 89
rect 202 88 203 89
rect 203 88 204 89
rect 204 88 205 89
rect 205 88 206 89
rect 206 88 207 89
rect 207 88 208 89
rect 208 88 209 89
rect 278 88 279 89
rect 279 88 280 89
rect 280 88 281 89
rect 281 88 282 89
rect 282 88 283 89
rect 283 88 284 89
rect 284 88 285 89
rect 285 88 286 89
rect 286 88 287 89
rect 287 88 288 89
rect 199 87 200 88
rect 200 87 201 88
rect 201 87 202 88
rect 202 87 203 88
rect 203 87 204 88
rect 204 87 205 88
rect 205 87 206 88
rect 206 87 207 88
rect 207 87 208 88
rect 208 87 209 88
rect 209 87 210 88
rect 277 87 278 88
rect 278 87 279 88
rect 279 87 280 88
rect 280 87 281 88
rect 281 87 282 88
rect 282 87 283 88
rect 283 87 284 88
rect 284 87 285 88
rect 285 87 286 88
rect 286 87 287 88
rect 200 86 201 87
rect 201 86 202 87
rect 202 86 203 87
rect 203 86 204 87
rect 204 86 205 87
rect 205 86 206 87
rect 206 86 207 87
rect 207 86 208 87
rect 208 86 209 87
rect 209 86 210 87
rect 210 86 211 87
rect 276 86 277 87
rect 277 86 278 87
rect 278 86 279 87
rect 279 86 280 87
rect 280 86 281 87
rect 281 86 282 87
rect 282 86 283 87
rect 283 86 284 87
rect 284 86 285 87
rect 285 86 286 87
rect 199 85 200 86
rect 200 85 201 86
rect 201 85 202 86
rect 202 85 203 86
rect 203 85 204 86
rect 204 85 205 86
rect 205 85 206 86
rect 206 85 207 86
rect 207 85 208 86
rect 208 85 209 86
rect 209 85 210 86
rect 210 85 211 86
rect 211 85 212 86
rect 275 85 276 86
rect 276 85 277 86
rect 277 85 278 86
rect 278 85 279 86
rect 279 85 280 86
rect 280 85 281 86
rect 281 85 282 86
rect 282 85 283 86
rect 283 85 284 86
rect 284 85 285 86
rect 199 84 200 85
rect 200 84 201 85
rect 201 84 202 85
rect 202 84 203 85
rect 203 84 204 85
rect 205 84 206 85
rect 206 84 207 85
rect 207 84 208 85
rect 208 84 209 85
rect 209 84 210 85
rect 210 84 211 85
rect 211 84 212 85
rect 275 84 276 85
rect 276 84 277 85
rect 277 84 278 85
rect 278 84 279 85
rect 279 84 280 85
rect 280 84 281 85
rect 281 84 282 85
rect 282 84 283 85
rect 283 84 284 85
rect 284 84 285 85
rect 199 83 200 84
rect 200 83 201 84
rect 201 83 202 84
rect 202 83 203 84
rect 203 83 204 84
rect 206 83 207 84
rect 207 83 208 84
rect 208 83 209 84
rect 209 83 210 84
rect 210 83 211 84
rect 211 83 212 84
rect 212 83 213 84
rect 274 83 275 84
rect 275 83 276 84
rect 276 83 277 84
rect 277 83 278 84
rect 278 83 279 84
rect 279 83 280 84
rect 280 83 281 84
rect 281 83 282 84
rect 282 83 283 84
rect 283 83 284 84
rect 199 82 200 83
rect 200 82 201 83
rect 201 82 202 83
rect 202 82 203 83
rect 203 82 204 83
rect 207 82 208 83
rect 208 82 209 83
rect 209 82 210 83
rect 210 82 211 83
rect 211 82 212 83
rect 212 82 213 83
rect 213 82 214 83
rect 273 82 274 83
rect 274 82 275 83
rect 275 82 276 83
rect 276 82 277 83
rect 277 82 278 83
rect 278 82 279 83
rect 279 82 280 83
rect 280 82 281 83
rect 281 82 282 83
rect 282 82 283 83
rect 198 81 199 82
rect 199 81 200 82
rect 200 81 201 82
rect 201 81 202 82
rect 202 81 203 82
rect 203 81 204 82
rect 208 81 209 82
rect 209 81 210 82
rect 210 81 211 82
rect 211 81 212 82
rect 212 81 213 82
rect 213 81 214 82
rect 214 81 215 82
rect 272 81 273 82
rect 273 81 274 82
rect 274 81 275 82
rect 275 81 276 82
rect 276 81 277 82
rect 277 81 278 82
rect 278 81 279 82
rect 279 81 280 82
rect 280 81 281 82
rect 281 81 282 82
rect 198 80 199 81
rect 199 80 200 81
rect 200 80 201 81
rect 201 80 202 81
rect 202 80 203 81
rect 203 80 204 81
rect 209 80 210 81
rect 210 80 211 81
rect 211 80 212 81
rect 212 80 213 81
rect 213 80 214 81
rect 214 80 215 81
rect 271 80 272 81
rect 272 80 273 81
rect 273 80 274 81
rect 274 80 275 81
rect 275 80 276 81
rect 276 80 277 81
rect 277 80 278 81
rect 278 80 279 81
rect 279 80 280 81
rect 280 80 281 81
rect 198 79 199 80
rect 199 79 200 80
rect 200 79 201 80
rect 201 79 202 80
rect 202 79 203 80
rect 203 79 204 80
rect 209 79 210 80
rect 210 79 211 80
rect 211 79 212 80
rect 212 79 213 80
rect 213 79 214 80
rect 214 79 215 80
rect 215 79 216 80
rect 270 79 271 80
rect 271 79 272 80
rect 272 79 273 80
rect 273 79 274 80
rect 274 79 275 80
rect 275 79 276 80
rect 276 79 277 80
rect 277 79 278 80
rect 278 79 279 80
rect 279 79 280 80
rect 198 78 199 79
rect 199 78 200 79
rect 200 78 201 79
rect 201 78 202 79
rect 202 78 203 79
rect 210 78 211 79
rect 211 78 212 79
rect 212 78 213 79
rect 213 78 214 79
rect 214 78 215 79
rect 215 78 216 79
rect 216 78 217 79
rect 269 78 270 79
rect 270 78 271 79
rect 271 78 272 79
rect 272 78 273 79
rect 273 78 274 79
rect 274 78 275 79
rect 275 78 276 79
rect 276 78 277 79
rect 277 78 278 79
rect 278 78 279 79
rect 197 77 198 78
rect 198 77 199 78
rect 199 77 200 78
rect 200 77 201 78
rect 201 77 202 78
rect 202 77 203 78
rect 211 77 212 78
rect 212 77 213 78
rect 213 77 214 78
rect 214 77 215 78
rect 215 77 216 78
rect 216 77 217 78
rect 268 77 269 78
rect 269 77 270 78
rect 270 77 271 78
rect 271 77 272 78
rect 272 77 273 78
rect 273 77 274 78
rect 274 77 275 78
rect 275 77 276 78
rect 276 77 277 78
rect 277 77 278 78
rect 278 77 279 78
rect 197 76 198 77
rect 198 76 199 77
rect 199 76 200 77
rect 200 76 201 77
rect 201 76 202 77
rect 202 76 203 77
rect 211 76 212 77
rect 212 76 213 77
rect 213 76 214 77
rect 214 76 215 77
rect 215 76 216 77
rect 216 76 217 77
rect 217 76 218 77
rect 268 76 269 77
rect 269 76 270 77
rect 270 76 271 77
rect 271 76 272 77
rect 272 76 273 77
rect 273 76 274 77
rect 274 76 275 77
rect 275 76 276 77
rect 276 76 277 77
rect 277 76 278 77
rect 196 75 197 76
rect 197 75 198 76
rect 198 75 199 76
rect 199 75 200 76
rect 200 75 201 76
rect 201 75 202 76
rect 202 75 203 76
rect 212 75 213 76
rect 213 75 214 76
rect 214 75 215 76
rect 215 75 216 76
rect 216 75 217 76
rect 217 75 218 76
rect 218 75 219 76
rect 267 75 268 76
rect 268 75 269 76
rect 269 75 270 76
rect 270 75 271 76
rect 271 75 272 76
rect 272 75 273 76
rect 273 75 274 76
rect 274 75 275 76
rect 275 75 276 76
rect 276 75 277 76
rect 196 74 197 75
rect 197 74 198 75
rect 198 74 199 75
rect 199 74 200 75
rect 200 74 201 75
rect 201 74 202 75
rect 213 74 214 75
rect 214 74 215 75
rect 215 74 216 75
rect 216 74 217 75
rect 217 74 218 75
rect 218 74 219 75
rect 266 74 267 75
rect 267 74 268 75
rect 268 74 269 75
rect 269 74 270 75
rect 270 74 271 75
rect 271 74 272 75
rect 272 74 273 75
rect 273 74 274 75
rect 274 74 275 75
rect 275 74 276 75
rect 196 73 197 74
rect 197 73 198 74
rect 198 73 199 74
rect 199 73 200 74
rect 200 73 201 74
rect 201 73 202 74
rect 213 73 214 74
rect 214 73 215 74
rect 215 73 216 74
rect 216 73 217 74
rect 217 73 218 74
rect 218 73 219 74
rect 219 73 220 74
rect 265 73 266 74
rect 266 73 267 74
rect 267 73 268 74
rect 268 73 269 74
rect 269 73 270 74
rect 270 73 271 74
rect 271 73 272 74
rect 272 73 273 74
rect 273 73 274 74
rect 274 73 275 74
rect 195 72 196 73
rect 196 72 197 73
rect 197 72 198 73
rect 198 72 199 73
rect 199 72 200 73
rect 200 72 201 73
rect 214 72 215 73
rect 215 72 216 73
rect 216 72 217 73
rect 217 72 218 73
rect 218 72 219 73
rect 219 72 220 73
rect 264 72 265 73
rect 265 72 266 73
rect 266 72 267 73
rect 267 72 268 73
rect 268 72 269 73
rect 269 72 270 73
rect 270 72 271 73
rect 271 72 272 73
rect 272 72 273 73
rect 273 72 274 73
rect 195 71 196 72
rect 196 71 197 72
rect 197 71 198 72
rect 198 71 199 72
rect 199 71 200 72
rect 200 71 201 72
rect 215 71 216 72
rect 216 71 217 72
rect 217 71 218 72
rect 218 71 219 72
rect 219 71 220 72
rect 220 71 221 72
rect 263 71 264 72
rect 264 71 265 72
rect 265 71 266 72
rect 266 71 267 72
rect 267 71 268 72
rect 268 71 269 72
rect 269 71 270 72
rect 270 71 271 72
rect 271 71 272 72
rect 272 71 273 72
rect 195 70 196 71
rect 196 70 197 71
rect 197 70 198 71
rect 198 70 199 71
rect 199 70 200 71
rect 200 70 201 71
rect 215 70 216 71
rect 216 70 217 71
rect 217 70 218 71
rect 218 70 219 71
rect 219 70 220 71
rect 220 70 221 71
rect 262 70 263 71
rect 263 70 264 71
rect 264 70 265 71
rect 265 70 266 71
rect 266 70 267 71
rect 267 70 268 71
rect 268 70 269 71
rect 269 70 270 71
rect 270 70 271 71
rect 271 70 272 71
rect 194 69 195 70
rect 195 69 196 70
rect 196 69 197 70
rect 197 69 198 70
rect 198 69 199 70
rect 199 69 200 70
rect 216 69 217 70
rect 217 69 218 70
rect 218 69 219 70
rect 219 69 220 70
rect 220 69 221 70
rect 221 69 222 70
rect 261 69 262 70
rect 262 69 263 70
rect 263 69 264 70
rect 264 69 265 70
rect 265 69 266 70
rect 266 69 267 70
rect 267 69 268 70
rect 268 69 269 70
rect 269 69 270 70
rect 270 69 271 70
rect 194 68 195 69
rect 195 68 196 69
rect 196 68 197 69
rect 197 68 198 69
rect 198 68 199 69
rect 199 68 200 69
rect 216 68 217 69
rect 217 68 218 69
rect 218 68 219 69
rect 219 68 220 69
rect 220 68 221 69
rect 221 68 222 69
rect 260 68 261 69
rect 261 68 262 69
rect 262 68 263 69
rect 263 68 264 69
rect 264 68 265 69
rect 265 68 266 69
rect 266 68 267 69
rect 267 68 268 69
rect 268 68 269 69
rect 269 68 270 69
rect 193 67 194 68
rect 194 67 195 68
rect 195 67 196 68
rect 196 67 197 68
rect 197 67 198 68
rect 198 67 199 68
rect 199 67 200 68
rect 217 67 218 68
rect 218 67 219 68
rect 219 67 220 68
rect 220 67 221 68
rect 221 67 222 68
rect 259 67 260 68
rect 260 67 261 68
rect 261 67 262 68
rect 262 67 263 68
rect 263 67 264 68
rect 264 67 265 68
rect 265 67 266 68
rect 266 67 267 68
rect 267 67 268 68
rect 268 67 269 68
rect 193 66 194 67
rect 194 66 195 67
rect 195 66 196 67
rect 196 66 197 67
rect 197 66 198 67
rect 198 66 199 67
rect 217 66 218 67
rect 218 66 219 67
rect 219 66 220 67
rect 220 66 221 67
rect 221 66 222 67
rect 222 66 223 67
rect 258 66 259 67
rect 259 66 260 67
rect 260 66 261 67
rect 261 66 262 67
rect 262 66 263 67
rect 263 66 264 67
rect 264 66 265 67
rect 265 66 266 67
rect 266 66 267 67
rect 267 66 268 67
rect 193 65 194 66
rect 194 65 195 66
rect 195 65 196 66
rect 196 65 197 66
rect 197 65 198 66
rect 198 65 199 66
rect 217 65 218 66
rect 218 65 219 66
rect 219 65 220 66
rect 220 65 221 66
rect 221 65 222 66
rect 222 65 223 66
rect 257 65 258 66
rect 258 65 259 66
rect 259 65 260 66
rect 260 65 261 66
rect 261 65 262 66
rect 262 65 263 66
rect 263 65 264 66
rect 264 65 265 66
rect 265 65 266 66
rect 266 65 267 66
rect 192 64 193 65
rect 193 64 194 65
rect 194 64 195 65
rect 195 64 196 65
rect 196 64 197 65
rect 197 64 198 65
rect 216 64 217 65
rect 217 64 218 65
rect 218 64 219 65
rect 219 64 220 65
rect 220 64 221 65
rect 221 64 222 65
rect 222 64 223 65
rect 256 64 257 65
rect 257 64 258 65
rect 258 64 259 65
rect 259 64 260 65
rect 260 64 261 65
rect 261 64 262 65
rect 262 64 263 65
rect 263 64 264 65
rect 264 64 265 65
rect 265 64 266 65
rect 192 63 193 64
rect 193 63 194 64
rect 194 63 195 64
rect 195 63 196 64
rect 196 63 197 64
rect 197 63 198 64
rect 214 63 215 64
rect 215 63 216 64
rect 216 63 217 64
rect 217 63 218 64
rect 218 63 219 64
rect 219 63 220 64
rect 220 63 221 64
rect 221 63 222 64
rect 222 63 223 64
rect 223 63 224 64
rect 255 63 256 64
rect 256 63 257 64
rect 257 63 258 64
rect 258 63 259 64
rect 259 63 260 64
rect 260 63 261 64
rect 261 63 262 64
rect 262 63 263 64
rect 263 63 264 64
rect 264 63 265 64
rect 191 62 192 63
rect 192 62 193 63
rect 193 62 194 63
rect 194 62 195 63
rect 195 62 196 63
rect 196 62 197 63
rect 197 62 198 63
rect 210 62 211 63
rect 211 62 212 63
rect 212 62 213 63
rect 213 62 214 63
rect 214 62 215 63
rect 215 62 216 63
rect 216 62 217 63
rect 217 62 218 63
rect 218 62 219 63
rect 219 62 220 63
rect 220 62 221 63
rect 221 62 222 63
rect 222 62 223 63
rect 223 62 224 63
rect 254 62 255 63
rect 255 62 256 63
rect 256 62 257 63
rect 257 62 258 63
rect 258 62 259 63
rect 259 62 260 63
rect 260 62 261 63
rect 261 62 262 63
rect 262 62 263 63
rect 263 62 264 63
rect 191 61 192 62
rect 192 61 193 62
rect 193 61 194 62
rect 194 61 195 62
rect 195 61 196 62
rect 196 61 197 62
rect 197 61 198 62
rect 198 61 199 62
rect 199 61 200 62
rect 200 61 201 62
rect 201 61 202 62
rect 202 61 203 62
rect 203 61 204 62
rect 204 61 205 62
rect 205 61 206 62
rect 206 61 207 62
rect 207 61 208 62
rect 208 61 209 62
rect 209 61 210 62
rect 210 61 211 62
rect 211 61 212 62
rect 212 61 213 62
rect 213 61 214 62
rect 214 61 215 62
rect 215 61 216 62
rect 216 61 217 62
rect 217 61 218 62
rect 218 61 219 62
rect 219 61 220 62
rect 220 61 221 62
rect 221 61 222 62
rect 222 61 223 62
rect 223 61 224 62
rect 253 61 254 62
rect 254 61 255 62
rect 255 61 256 62
rect 256 61 257 62
rect 257 61 258 62
rect 258 61 259 62
rect 259 61 260 62
rect 260 61 261 62
rect 261 61 262 62
rect 262 61 263 62
rect 191 60 192 61
rect 192 60 193 61
rect 193 60 194 61
rect 194 60 195 61
rect 195 60 196 61
rect 196 60 197 61
rect 197 60 198 61
rect 198 60 199 61
rect 199 60 200 61
rect 200 60 201 61
rect 201 60 202 61
rect 202 60 203 61
rect 203 60 204 61
rect 204 60 205 61
rect 205 60 206 61
rect 206 60 207 61
rect 207 60 208 61
rect 208 60 209 61
rect 209 60 210 61
rect 210 60 211 61
rect 211 60 212 61
rect 212 60 213 61
rect 213 60 214 61
rect 214 60 215 61
rect 215 60 216 61
rect 216 60 217 61
rect 217 60 218 61
rect 218 60 219 61
rect 219 60 220 61
rect 220 60 221 61
rect 221 60 222 61
rect 222 60 223 61
rect 223 60 224 61
rect 224 60 225 61
rect 252 60 253 61
rect 253 60 254 61
rect 254 60 255 61
rect 255 60 256 61
rect 256 60 257 61
rect 257 60 258 61
rect 258 60 259 61
rect 259 60 260 61
rect 260 60 261 61
rect 261 60 262 61
rect 190 59 191 60
rect 191 59 192 60
rect 192 59 193 60
rect 193 59 194 60
rect 194 59 195 60
rect 195 59 196 60
rect 196 59 197 60
rect 197 59 198 60
rect 198 59 199 60
rect 199 59 200 60
rect 200 59 201 60
rect 201 59 202 60
rect 202 59 203 60
rect 203 59 204 60
rect 204 59 205 60
rect 205 59 206 60
rect 206 59 207 60
rect 207 59 208 60
rect 208 59 209 60
rect 209 59 210 60
rect 210 59 211 60
rect 211 59 212 60
rect 212 59 213 60
rect 213 59 214 60
rect 214 59 215 60
rect 215 59 216 60
rect 216 59 217 60
rect 217 59 218 60
rect 218 59 219 60
rect 219 59 220 60
rect 220 59 221 60
rect 221 59 222 60
rect 222 59 223 60
rect 223 59 224 60
rect 224 59 225 60
rect 251 59 252 60
rect 252 59 253 60
rect 253 59 254 60
rect 254 59 255 60
rect 255 59 256 60
rect 256 59 257 60
rect 257 59 258 60
rect 258 59 259 60
rect 259 59 260 60
rect 260 59 261 60
rect 191 58 192 59
rect 192 58 193 59
rect 193 58 194 59
rect 194 58 195 59
rect 195 58 196 59
rect 196 58 197 59
rect 197 58 198 59
rect 198 58 199 59
rect 199 58 200 59
rect 200 58 201 59
rect 201 58 202 59
rect 202 58 203 59
rect 203 58 204 59
rect 204 58 205 59
rect 205 58 206 59
rect 206 58 207 59
rect 207 58 208 59
rect 208 58 209 59
rect 209 58 210 59
rect 210 58 211 59
rect 211 58 212 59
rect 212 58 213 59
rect 213 58 214 59
rect 214 58 215 59
rect 217 58 218 59
rect 218 58 219 59
rect 219 58 220 59
rect 220 58 221 59
rect 221 58 222 59
rect 222 58 223 59
rect 223 58 224 59
rect 224 58 225 59
rect 250 58 251 59
rect 251 58 252 59
rect 252 58 253 59
rect 253 58 254 59
rect 254 58 255 59
rect 255 58 256 59
rect 256 58 257 59
rect 257 58 258 59
rect 258 58 259 59
rect 259 58 260 59
rect 191 57 192 58
rect 192 57 193 58
rect 193 57 194 58
rect 194 57 195 58
rect 195 57 196 58
rect 196 57 197 58
rect 197 57 198 58
rect 198 57 199 58
rect 199 57 200 58
rect 200 57 201 58
rect 201 57 202 58
rect 202 57 203 58
rect 203 57 204 58
rect 204 57 205 58
rect 205 57 206 58
rect 206 57 207 58
rect 207 57 208 58
rect 208 57 209 58
rect 209 57 210 58
rect 210 57 211 58
rect 211 57 212 58
rect 212 57 213 58
rect 217 57 218 58
rect 218 57 219 58
rect 219 57 220 58
rect 220 57 221 58
rect 221 57 222 58
rect 222 57 223 58
rect 223 57 224 58
rect 224 57 225 58
rect 249 57 250 58
rect 250 57 251 58
rect 251 57 252 58
rect 252 57 253 58
rect 253 57 254 58
rect 254 57 255 58
rect 255 57 256 58
rect 256 57 257 58
rect 257 57 258 58
rect 258 57 259 58
rect 191 56 192 57
rect 192 56 193 57
rect 193 56 194 57
rect 194 56 195 57
rect 195 56 196 57
rect 196 56 197 57
rect 197 56 198 57
rect 198 56 199 57
rect 199 56 200 57
rect 200 56 201 57
rect 201 56 202 57
rect 202 56 203 57
rect 203 56 204 57
rect 204 56 205 57
rect 205 56 206 57
rect 206 56 207 57
rect 207 56 208 57
rect 208 56 209 57
rect 209 56 210 57
rect 217 56 218 57
rect 218 56 219 57
rect 219 56 220 57
rect 220 56 221 57
rect 221 56 222 57
rect 222 56 223 57
rect 223 56 224 57
rect 224 56 225 57
rect 248 56 249 57
rect 249 56 250 57
rect 250 56 251 57
rect 251 56 252 57
rect 252 56 253 57
rect 253 56 254 57
rect 254 56 255 57
rect 255 56 256 57
rect 256 56 257 57
rect 257 56 258 57
rect 193 55 194 56
rect 194 55 195 56
rect 195 55 196 56
rect 196 55 197 56
rect 197 55 198 56
rect 198 55 199 56
rect 199 55 200 56
rect 200 55 201 56
rect 201 55 202 56
rect 202 55 203 56
rect 203 55 204 56
rect 204 55 205 56
rect 205 55 206 56
rect 206 55 207 56
rect 217 55 218 56
rect 218 55 219 56
rect 219 55 220 56
rect 220 55 221 56
rect 221 55 222 56
rect 222 55 223 56
rect 223 55 224 56
rect 224 55 225 56
rect 247 55 248 56
rect 248 55 249 56
rect 249 55 250 56
rect 250 55 251 56
rect 251 55 252 56
rect 252 55 253 56
rect 253 55 254 56
rect 254 55 255 56
rect 255 55 256 56
rect 256 55 257 56
rect 198 54 199 55
rect 199 54 200 55
rect 217 54 218 55
rect 218 54 219 55
rect 219 54 220 55
rect 220 54 221 55
rect 221 54 222 55
rect 222 54 223 55
rect 223 54 224 55
rect 224 54 225 55
rect 246 54 247 55
rect 247 54 248 55
rect 248 54 249 55
rect 249 54 250 55
rect 250 54 251 55
rect 251 54 252 55
rect 252 54 253 55
rect 253 54 254 55
rect 254 54 255 55
rect 255 54 256 55
rect 218 53 219 54
rect 219 53 220 54
rect 220 53 221 54
rect 221 53 222 54
rect 222 53 223 54
rect 223 53 224 54
rect 224 53 225 54
rect 225 53 226 54
rect 245 53 246 54
rect 246 53 247 54
rect 247 53 248 54
rect 248 53 249 54
rect 249 53 250 54
rect 250 53 251 54
rect 251 53 252 54
rect 252 53 253 54
rect 253 53 254 54
rect 254 53 255 54
rect 218 52 219 53
rect 219 52 220 53
rect 220 52 221 53
rect 221 52 222 53
rect 222 52 223 53
rect 223 52 224 53
rect 224 52 225 53
rect 225 52 226 53
rect 244 52 245 53
rect 245 52 246 53
rect 246 52 247 53
rect 247 52 248 53
rect 248 52 249 53
rect 249 52 250 53
rect 250 52 251 53
rect 251 52 252 53
rect 252 52 253 53
rect 253 52 254 53
rect 218 51 219 52
rect 219 51 220 52
rect 220 51 221 52
rect 221 51 222 52
rect 222 51 223 52
rect 223 51 224 52
rect 224 51 225 52
rect 225 51 226 52
rect 243 51 244 52
rect 244 51 245 52
rect 245 51 246 52
rect 246 51 247 52
rect 247 51 248 52
rect 248 51 249 52
rect 249 51 250 52
rect 250 51 251 52
rect 251 51 252 52
rect 252 51 253 52
rect 218 50 219 51
rect 219 50 220 51
rect 220 50 221 51
rect 221 50 222 51
rect 222 50 223 51
rect 223 50 224 51
rect 224 50 225 51
rect 225 50 226 51
rect 242 50 243 51
rect 243 50 244 51
rect 244 50 245 51
rect 245 50 246 51
rect 246 50 247 51
rect 247 50 248 51
rect 248 50 249 51
rect 249 50 250 51
rect 250 50 251 51
rect 251 50 252 51
rect 218 49 219 50
rect 219 49 220 50
rect 220 49 221 50
rect 221 49 222 50
rect 222 49 223 50
rect 223 49 224 50
rect 224 49 225 50
rect 225 49 226 50
rect 241 49 242 50
rect 242 49 243 50
rect 243 49 244 50
rect 244 49 245 50
rect 245 49 246 50
rect 246 49 247 50
rect 247 49 248 50
rect 248 49 249 50
rect 249 49 250 50
rect 250 49 251 50
rect 218 48 219 49
rect 219 48 220 49
rect 220 48 221 49
rect 221 48 222 49
rect 222 48 223 49
rect 223 48 224 49
rect 224 48 225 49
rect 225 48 226 49
rect 240 48 241 49
rect 241 48 242 49
rect 242 48 243 49
rect 243 48 244 49
rect 244 48 245 49
rect 245 48 246 49
rect 246 48 247 49
rect 247 48 248 49
rect 248 48 249 49
rect 249 48 250 49
rect 218 47 219 48
rect 219 47 220 48
rect 220 47 221 48
rect 221 47 222 48
rect 222 47 223 48
rect 223 47 224 48
rect 224 47 225 48
rect 225 47 226 48
rect 239 47 240 48
rect 240 47 241 48
rect 241 47 242 48
rect 242 47 243 48
rect 243 47 244 48
rect 244 47 245 48
rect 245 47 246 48
rect 246 47 247 48
rect 247 47 248 48
rect 248 47 249 48
rect 219 46 220 47
rect 220 46 221 47
rect 221 46 222 47
rect 222 46 223 47
rect 223 46 224 47
rect 224 46 225 47
rect 225 46 226 47
rect 238 46 239 47
rect 239 46 240 47
rect 240 46 241 47
rect 241 46 242 47
rect 242 46 243 47
rect 243 46 244 47
rect 244 46 245 47
rect 245 46 246 47
rect 246 46 247 47
rect 247 46 248 47
rect 219 45 220 46
rect 220 45 221 46
rect 221 45 222 46
rect 222 45 223 46
rect 223 45 224 46
rect 224 45 225 46
rect 225 45 226 46
rect 237 45 238 46
rect 238 45 239 46
rect 239 45 240 46
rect 240 45 241 46
rect 241 45 242 46
rect 242 45 243 46
rect 243 45 244 46
rect 244 45 245 46
rect 245 45 246 46
rect 246 45 247 46
rect 219 44 220 45
rect 220 44 221 45
rect 221 44 222 45
rect 222 44 223 45
rect 223 44 224 45
rect 224 44 225 45
rect 225 44 226 45
rect 236 44 237 45
rect 237 44 238 45
rect 238 44 239 45
rect 239 44 240 45
rect 240 44 241 45
rect 241 44 242 45
rect 242 44 243 45
rect 243 44 244 45
rect 244 44 245 45
rect 245 44 246 45
rect 219 43 220 44
rect 220 43 221 44
rect 221 43 222 44
rect 222 43 223 44
rect 223 43 224 44
rect 224 43 225 44
rect 225 43 226 44
rect 235 43 236 44
rect 236 43 237 44
rect 237 43 238 44
rect 238 43 239 44
rect 239 43 240 44
rect 240 43 241 44
rect 241 43 242 44
rect 242 43 243 44
rect 243 43 244 44
rect 244 43 245 44
rect 219 42 220 43
rect 220 42 221 43
rect 221 42 222 43
rect 222 42 223 43
rect 223 42 224 43
rect 224 42 225 43
rect 225 42 226 43
rect 233 42 234 43
rect 234 42 235 43
rect 235 42 236 43
rect 236 42 237 43
rect 237 42 238 43
rect 238 42 239 43
rect 239 42 240 43
rect 240 42 241 43
rect 241 42 242 43
rect 242 42 243 43
rect 243 42 244 43
rect 219 41 220 42
rect 220 41 221 42
rect 221 41 222 42
rect 222 41 223 42
rect 223 41 224 42
rect 224 41 225 42
rect 225 41 226 42
rect 232 41 233 42
rect 233 41 234 42
rect 234 41 235 42
rect 235 41 236 42
rect 236 41 237 42
rect 237 41 238 42
rect 238 41 239 42
rect 239 41 240 42
rect 240 41 241 42
rect 241 41 242 42
rect 242 41 243 42
rect 219 40 220 41
rect 220 40 221 41
rect 221 40 222 41
rect 222 40 223 41
rect 223 40 224 41
rect 224 40 225 41
rect 225 40 226 41
rect 231 40 232 41
rect 232 40 233 41
rect 233 40 234 41
rect 234 40 235 41
rect 235 40 236 41
rect 236 40 237 41
rect 237 40 238 41
rect 238 40 239 41
rect 239 40 240 41
rect 240 40 241 41
rect 241 40 242 41
rect 219 39 220 40
rect 220 39 221 40
rect 221 39 222 40
rect 222 39 223 40
rect 223 39 224 40
rect 224 39 225 40
rect 225 39 226 40
rect 230 39 231 40
rect 231 39 232 40
rect 232 39 233 40
rect 233 39 234 40
rect 234 39 235 40
rect 235 39 236 40
rect 236 39 237 40
rect 237 39 238 40
rect 238 39 239 40
rect 239 39 240 40
rect 240 39 241 40
rect 219 38 220 39
rect 220 38 221 39
rect 221 38 222 39
rect 222 38 223 39
rect 223 38 224 39
rect 224 38 225 39
rect 225 38 226 39
rect 226 38 227 39
rect 227 38 228 39
rect 228 38 229 39
rect 229 38 230 39
rect 230 38 231 39
rect 231 38 232 39
rect 232 38 233 39
rect 233 38 234 39
rect 234 38 235 39
rect 235 38 236 39
rect 236 38 237 39
rect 237 38 238 39
rect 238 38 239 39
rect 219 37 220 38
rect 220 37 221 38
rect 221 37 222 38
rect 222 37 223 38
rect 223 37 224 38
rect 224 37 225 38
rect 225 37 226 38
rect 226 37 227 38
rect 227 37 228 38
rect 228 37 229 38
rect 229 37 230 38
rect 230 37 231 38
rect 231 37 232 38
rect 232 37 233 38
rect 233 37 234 38
rect 234 37 235 38
rect 235 37 236 38
rect 236 37 237 38
rect 237 37 238 38
rect 220 36 221 37
rect 221 36 222 37
rect 222 36 223 37
rect 223 36 224 37
rect 224 36 225 37
rect 225 36 226 37
rect 226 36 227 37
rect 227 36 228 37
rect 228 36 229 37
rect 229 36 230 37
rect 230 36 231 37
rect 231 36 232 37
rect 232 36 233 37
rect 233 36 234 37
rect 234 36 235 37
rect 235 36 236 37
rect 236 36 237 37
rect 220 35 221 36
rect 221 35 222 36
rect 222 35 223 36
rect 223 35 224 36
rect 224 35 225 36
rect 225 35 226 36
rect 226 35 227 36
rect 227 35 228 36
rect 228 35 229 36
rect 229 35 230 36
rect 230 35 231 36
rect 231 35 232 36
rect 232 35 233 36
rect 233 35 234 36
rect 234 35 235 36
rect 235 35 236 36
rect 220 34 221 35
rect 221 34 222 35
rect 222 34 223 35
rect 223 34 224 35
rect 224 34 225 35
rect 225 34 226 35
rect 226 34 227 35
rect 227 34 228 35
rect 228 34 229 35
rect 229 34 230 35
rect 230 34 231 35
rect 231 34 232 35
rect 232 34 233 35
rect 233 34 234 35
rect 234 34 235 35
rect 221 33 222 34
rect 222 33 223 34
rect 223 33 224 34
rect 224 33 225 34
rect 225 33 226 34
rect 226 33 227 34
rect 227 33 228 34
rect 228 33 229 34
rect 229 33 230 34
rect 230 33 231 34
rect 231 33 232 34
rect 232 33 233 34
rect 233 33 234 34
rect 221 32 222 33
rect 222 32 223 33
rect 223 32 224 33
rect 224 32 225 33
rect 225 32 226 33
rect 226 32 227 33
rect 227 32 228 33
rect 228 32 229 33
rect 229 32 230 33
rect 230 32 231 33
rect 231 32 232 33
rect 232 32 233 33
rect 223 31 224 32
rect 224 31 225 32
rect 225 31 226 32
rect 226 31 227 32
rect 227 31 228 32
rect 228 31 229 32
rect 229 31 230 32
rect 230 31 231 32
rect 231 31 232 32
rect 227 30 228 31
rect 228 30 229 31
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1606864417
<< checkpaint >>
rect -1209 -1243 2569 2131
<< nwell >>
rect -9 485 1435 897
<< nmos >>
rect 80 115 110 219
rect 166 115 196 219
rect 252 115 282 219
rect 338 115 368 219
rect 410 115 440 219
rect 496 115 526 219
rect 582 115 612 219
rect 668 115 698 219
rect 754 115 784 219
rect 840 115 870 219
rect 922 115 952 219
rect 1004 115 1034 219
rect 1102 115 1132 219
rect 1292 115 1322 219
<< pmos >>
rect 80 521 110 773
rect 166 521 196 773
rect 252 521 282 773
rect 338 521 368 773
rect 410 521 440 773
rect 496 521 526 773
rect 582 521 612 773
rect 668 521 698 773
rect 754 521 784 773
rect 840 521 870 773
rect 922 521 952 773
rect 1004 521 1034 773
rect 1102 521 1132 773
rect 1292 521 1322 773
<< ndiff >>
rect 27 171 80 219
rect 27 131 35 171
rect 69 131 80 171
rect 27 115 80 131
rect 110 165 166 219
rect 110 131 121 165
rect 155 131 166 165
rect 110 115 166 131
rect 196 171 252 219
rect 196 131 207 171
rect 241 131 252 171
rect 196 115 252 131
rect 282 171 338 219
rect 282 131 293 171
rect 327 131 338 171
rect 282 115 338 131
rect 368 115 410 219
rect 440 171 496 219
rect 440 131 451 171
rect 485 131 496 171
rect 440 115 496 131
rect 526 171 582 219
rect 526 131 537 171
rect 571 131 582 171
rect 526 115 582 131
rect 612 157 668 219
rect 612 123 623 157
rect 657 123 668 157
rect 612 115 668 123
rect 698 171 754 219
rect 698 131 709 171
rect 743 131 754 171
rect 698 115 754 131
rect 784 165 840 219
rect 784 131 795 165
rect 829 131 840 165
rect 784 115 840 131
rect 870 115 922 219
rect 952 115 1004 219
rect 1034 171 1102 219
rect 1034 131 1045 171
rect 1079 131 1102 171
rect 1034 115 1102 131
rect 1132 171 1185 219
rect 1132 131 1143 171
rect 1177 131 1185 171
rect 1132 115 1185 131
rect 1239 165 1292 219
rect 1239 131 1247 165
rect 1281 131 1292 165
rect 1239 115 1292 131
rect 1322 171 1375 219
rect 1322 131 1333 171
rect 1367 131 1375 171
rect 1322 115 1375 131
<< pdiff >>
rect 27 757 80 773
rect 27 629 35 757
rect 69 629 80 757
rect 27 521 80 629
rect 110 757 166 773
rect 110 697 121 757
rect 155 697 166 757
rect 110 521 166 697
rect 196 757 252 773
rect 196 629 207 757
rect 241 629 252 757
rect 196 521 252 629
rect 282 757 338 773
rect 282 629 293 757
rect 327 629 338 757
rect 282 521 338 629
rect 368 521 410 773
rect 440 757 496 773
rect 440 629 451 757
rect 485 629 496 757
rect 440 521 496 629
rect 526 757 582 773
rect 526 629 537 757
rect 571 629 582 757
rect 526 521 582 629
rect 612 757 668 773
rect 612 723 623 757
rect 657 723 668 757
rect 612 521 668 723
rect 698 757 754 773
rect 698 663 709 757
rect 743 663 754 757
rect 698 521 754 663
rect 784 757 840 773
rect 784 629 795 757
rect 829 629 840 757
rect 784 521 840 629
rect 870 521 922 773
rect 952 521 1004 773
rect 1034 757 1102 773
rect 1034 697 1045 757
rect 1079 697 1102 757
rect 1034 521 1102 697
rect 1132 757 1185 773
rect 1132 629 1143 757
rect 1177 629 1185 757
rect 1132 521 1185 629
rect 1239 757 1292 773
rect 1239 561 1247 757
rect 1281 561 1292 757
rect 1239 521 1292 561
rect 1322 757 1375 773
rect 1322 561 1333 757
rect 1367 561 1375 757
rect 1322 521 1375 561
<< ndiffc >>
rect 35 131 69 171
rect 121 131 155 165
rect 207 131 241 171
rect 293 131 327 171
rect 451 131 485 171
rect 537 131 571 171
rect 623 123 657 157
rect 709 131 743 171
rect 795 131 829 165
rect 1045 131 1079 171
rect 1143 131 1177 171
rect 1247 131 1281 165
rect 1333 131 1367 171
<< pdiffc >>
rect 35 629 69 757
rect 121 697 155 757
rect 207 629 241 757
rect 293 629 327 757
rect 451 629 485 757
rect 537 629 571 757
rect 623 723 657 757
rect 709 663 743 757
rect 795 629 829 757
rect 1045 697 1079 757
rect 1143 629 1177 757
rect 1247 561 1281 757
rect 1333 561 1367 757
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
rect 571 27 595 61
rect 629 27 653 61
rect 707 27 731 61
rect 765 27 789 61
rect 843 27 867 61
rect 901 27 925 61
rect 979 27 1003 61
rect 1037 27 1061 61
rect 1115 27 1139 61
rect 1173 27 1197 61
rect 1251 27 1275 61
rect 1309 27 1333 61
<< nsubdiff >>
rect 27 827 51 861
rect 85 827 109 861
rect 163 827 187 861
rect 221 827 245 861
rect 299 827 323 861
rect 357 827 381 861
rect 435 827 459 861
rect 493 827 517 861
rect 571 827 595 861
rect 629 827 653 861
rect 707 827 731 861
rect 765 827 789 861
rect 843 827 867 861
rect 901 827 925 861
rect 979 827 1003 861
rect 1037 827 1061 861
rect 1115 827 1139 861
rect 1173 827 1197 861
rect 1251 827 1275 861
rect 1309 827 1333 861
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
rect 595 27 629 61
rect 731 27 765 61
rect 867 27 901 61
rect 1003 27 1037 61
rect 1139 27 1173 61
rect 1275 27 1309 61
<< nsubdiffcont >>
rect 51 827 85 861
rect 187 827 221 861
rect 323 827 357 861
rect 459 827 493 861
rect 595 827 629 861
rect 731 827 765 861
rect 867 827 901 861
rect 1003 827 1037 861
rect 1139 827 1173 861
rect 1275 827 1309 861
<< poly >>
rect 80 773 110 799
rect 166 773 196 799
rect 252 773 282 801
rect 338 773 368 801
rect 410 773 440 799
rect 496 773 526 799
rect 582 773 612 801
rect 668 773 698 801
rect 754 773 784 801
rect 840 773 870 801
rect 922 773 952 801
rect 1004 773 1034 801
rect 1102 773 1132 801
rect 1292 773 1322 801
rect 80 381 110 521
rect 166 489 196 521
rect 152 473 206 489
rect 152 439 162 473
rect 196 439 206 473
rect 152 423 206 439
rect 70 365 124 381
rect 70 331 80 365
rect 114 331 124 365
rect 70 315 124 331
rect 80 219 110 315
rect 166 219 196 423
rect 252 381 282 521
rect 338 423 368 521
rect 410 496 440 521
rect 496 496 526 521
rect 410 466 526 496
rect 338 407 430 423
rect 238 365 292 381
rect 238 331 248 365
rect 282 331 292 365
rect 238 315 292 331
rect 338 373 386 407
rect 420 373 430 407
rect 338 357 430 373
rect 472 363 502 466
rect 582 364 612 521
rect 668 455 698 521
rect 656 439 710 455
rect 656 405 666 439
rect 700 405 710 439
rect 656 389 710 405
rect 252 219 282 315
rect 338 219 368 357
rect 472 347 526 363
rect 472 313 482 347
rect 516 313 526 347
rect 472 271 526 313
rect 568 348 622 364
rect 568 314 578 348
rect 612 314 622 348
rect 568 298 622 314
rect 410 241 526 271
rect 410 219 440 241
rect 496 219 526 241
rect 582 219 612 298
rect 668 219 698 389
rect 754 324 784 521
rect 840 460 870 521
rect 826 444 880 460
rect 826 410 836 444
rect 870 410 880 444
rect 826 394 880 410
rect 922 417 952 521
rect 1004 489 1034 521
rect 1004 459 1048 489
rect 1102 488 1132 521
rect 922 401 976 417
rect 742 308 796 324
rect 742 274 752 308
rect 786 274 796 308
rect 742 258 796 274
rect 754 219 784 258
rect 840 219 870 394
rect 922 367 932 401
rect 966 367 976 401
rect 922 351 976 367
rect 922 219 952 351
rect 1018 307 1048 459
rect 1090 472 1144 488
rect 1292 485 1322 521
rect 1090 438 1100 472
rect 1134 438 1144 472
rect 1090 422 1144 438
rect 1255 469 1322 485
rect 1255 435 1265 469
rect 1299 435 1322 469
rect 1004 291 1058 307
rect 1004 257 1014 291
rect 1048 257 1058 291
rect 1004 241 1058 257
rect 1004 219 1034 241
rect 1102 219 1132 422
rect 1255 419 1322 435
rect 1292 219 1322 419
rect 80 81 110 115
rect 166 82 196 115
rect 252 82 282 115
rect 338 82 368 115
rect 410 82 440 115
rect 496 82 526 115
rect 582 82 612 115
rect 668 82 698 115
rect 754 82 784 115
rect 840 82 870 115
rect 922 82 952 115
rect 1004 82 1034 115
rect 1102 80 1132 115
rect 1292 80 1322 115
<< polycont >>
rect 162 439 196 473
rect 80 331 114 365
rect 248 331 282 365
rect 386 373 420 407
rect 666 405 700 439
rect 482 313 516 347
rect 578 314 612 348
rect 836 410 870 444
rect 752 274 786 308
rect 932 367 966 401
rect 1100 438 1134 472
rect 1265 435 1299 469
rect 1014 257 1048 291
<< locali >>
rect 0 867 1408 888
rect 0 827 51 867
rect 85 827 187 867
rect 221 827 323 867
rect 357 827 459 867
rect 493 827 595 867
rect 629 827 731 867
rect 765 827 867 867
rect 901 827 1003 867
rect 1037 827 1139 867
rect 1173 827 1275 867
rect 1309 827 1408 867
rect 35 757 69 773
rect 121 757 155 827
rect 121 681 155 697
rect 207 757 241 773
rect 35 613 69 629
rect 207 613 241 629
rect 35 579 241 613
rect 293 757 327 773
rect 293 546 327 629
rect 451 757 485 827
rect 451 613 485 629
rect 537 757 571 773
rect 623 757 657 827
rect 623 707 657 723
rect 709 757 743 773
rect 571 629 743 663
rect 795 757 829 773
rect 1045 757 1079 827
rect 1045 681 1079 697
rect 1143 757 1177 773
rect 537 613 571 629
rect 795 588 829 629
rect 1143 588 1177 629
rect 752 554 1100 588
rect 752 553 812 554
rect 293 509 350 546
rect 80 473 114 479
rect 80 439 162 473
rect 196 439 212 473
rect 248 365 282 405
rect 64 331 80 365
rect 114 331 130 365
rect 248 315 282 331
rect 316 291 350 509
rect 386 479 444 513
rect 386 407 420 479
rect 386 357 420 373
rect 578 348 612 479
rect 752 510 787 553
rect 650 405 666 439
rect 700 405 716 439
rect 466 313 482 347
rect 516 313 532 347
rect 752 376 786 510
rect 836 444 870 479
rect 1066 488 1100 554
rect 1247 757 1281 827
rect 1177 554 1202 571
rect 1143 537 1202 554
rect 1247 545 1281 561
rect 1333 757 1367 773
rect 1066 472 1134 488
rect 820 410 836 444
rect 870 410 886 444
rect 1066 441 1100 472
rect 1089 438 1100 441
rect 1100 422 1134 438
rect 932 401 966 405
rect 752 342 879 376
rect 932 351 966 367
rect 1168 365 1202 537
rect 1333 513 1367 561
rect 578 298 612 314
rect 736 274 752 308
rect 786 291 810 308
rect 35 215 241 249
rect 35 189 70 215
rect 35 171 69 189
rect 35 115 69 131
rect 121 165 155 181
rect 121 61 155 131
rect 207 171 241 215
rect 207 114 241 131
rect 293 223 350 257
rect 293 171 327 223
rect 537 206 743 240
rect 293 114 327 131
rect 451 171 485 187
rect 451 61 485 131
rect 537 171 571 206
rect 709 171 743 206
rect 845 190 879 342
rect 1014 291 1048 331
rect 1143 331 1202 365
rect 1265 469 1299 485
rect 998 257 1014 291
rect 1048 257 1064 291
rect 1014 256 1048 257
rect 537 114 571 131
rect 607 123 623 157
rect 657 123 673 157
rect 623 61 657 123
rect 709 114 743 131
rect 795 165 879 190
rect 829 156 879 165
rect 1045 171 1079 187
rect 795 114 829 131
rect 1045 61 1079 131
rect 1143 171 1177 331
rect 1265 291 1299 435
rect 1245 257 1299 291
rect 1143 115 1177 131
rect 1247 165 1281 181
rect 1247 61 1281 131
rect 1333 171 1367 479
rect 1333 115 1367 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 595 61
rect 629 21 731 61
rect 765 21 867 61
rect 901 21 1003 61
rect 1037 21 1139 61
rect 1173 21 1275 61
rect 1309 21 1408 61
rect 0 0 1408 21
<< viali >>
rect 51 861 85 867
rect 51 833 85 861
rect 187 861 221 867
rect 187 833 221 861
rect 323 861 357 867
rect 323 833 357 861
rect 459 861 493 867
rect 459 833 493 861
rect 595 861 629 867
rect 595 833 629 861
rect 731 861 765 867
rect 731 833 765 861
rect 867 861 901 867
rect 867 833 901 861
rect 1003 861 1037 867
rect 1003 833 1037 861
rect 1139 861 1173 867
rect 1139 833 1173 861
rect 1275 861 1309 867
rect 1275 833 1309 861
rect 80 479 114 513
rect 248 405 282 439
rect 80 331 114 365
rect 444 479 478 513
rect 578 479 612 513
rect 482 347 516 365
rect 666 405 700 439
rect 482 331 516 347
rect 836 479 870 513
rect 1143 554 1177 588
rect 932 405 966 439
rect 316 257 350 291
rect 777 274 786 291
rect 786 274 811 291
rect 777 257 811 274
rect 1014 331 1048 365
rect 1211 257 1245 291
rect 1333 479 1367 513
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
rect 595 27 629 55
rect 595 21 629 27
rect 731 27 765 55
rect 731 21 765 27
rect 867 27 901 55
rect 867 21 901 27
rect 1003 27 1037 55
rect 1003 21 1037 27
rect 1139 27 1173 55
rect 1139 21 1173 27
rect 1275 27 1309 55
rect 1275 21 1309 27
<< metal1 >>
rect 0 867 1408 888
rect 0 833 51 867
rect 85 833 187 867
rect 221 833 323 867
rect 357 833 459 867
rect 493 833 595 867
rect 629 833 731 867
rect 765 833 867 867
rect 901 833 1003 867
rect 1037 833 1139 867
rect 1173 833 1275 867
rect 1309 833 1408 867
rect 0 827 1408 833
rect 1131 588 1189 594
rect 1109 554 1143 588
rect 1177 554 1189 588
rect 1131 548 1189 554
rect 68 513 126 519
rect 432 513 490 519
rect 566 513 624 519
rect 824 513 882 520
rect 1321 513 1379 519
rect 68 479 80 513
rect 114 479 444 513
rect 478 479 578 513
rect 612 479 836 513
rect 870 479 882 513
rect 1299 479 1333 513
rect 1367 479 1379 513
rect 68 473 126 479
rect 432 473 490 479
rect 566 473 624 479
rect 824 472 882 479
rect 1321 473 1379 479
rect 236 439 296 445
rect 650 439 717 445
rect 920 439 978 445
rect 236 405 248 439
rect 282 405 666 439
rect 700 405 932 439
rect 966 405 978 439
rect 236 399 296 405
rect 650 399 717 405
rect 920 399 978 405
rect 68 365 126 371
rect 470 365 528 371
rect 1002 365 1060 371
rect 68 331 80 365
rect 114 331 482 365
rect 516 331 1014 365
rect 1048 331 1060 365
rect 68 325 126 331
rect 470 325 528 331
rect 1002 325 1060 331
rect 304 291 362 297
rect 771 291 820 297
rect 1199 291 1257 297
rect 304 257 316 291
rect 350 257 777 291
rect 811 257 1211 291
rect 1245 257 1257 291
rect 304 251 362 257
rect 771 251 820 257
rect 1199 251 1257 257
rect 0 55 1408 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 595 55
rect 629 21 731 55
rect 765 21 867 55
rect 901 21 1003 55
rect 1037 21 1139 55
rect 1173 21 1275 55
rect 1309 21 1408 55
rect 0 0 1408 21
<< labels >>
rlabel viali 1160 571 1160 571 1 S
port 5 n
rlabel viali 1350 496 1350 496 1 CO
port 6 n
rlabel metal1 129 496 129 496 1 B
rlabel viali 265 422 265 422 1 CI
rlabel viali 97 348 97 348 1 A
port 1 n
rlabel viali 1228 274 1228 274 1 CON
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 840 68 840 1 vdd
<< end >>

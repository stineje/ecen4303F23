* FILE: top.sp

********************** begin header *****************************

* SPICE Header file for SKY130 process (sky130)

.OPTIONS post NOMOD probe measout captab 

**################################################
* Only Typical/Typical spice models included
.include '/programs/micromagic/mmi_local/ami05.mod'
**################################################

.param ln_min   =  0.15u
.param lp_min   =  0.15u

.PARAM vddp=3.30	$ VDD voltage

VDD vdd 0 DC vddp 

.TEMP 25
.TRAN 5p 10n

*********************** end header ******************************

* SPICE netlist for "top" generated by MMI_SUE5.6.41 on Thu Nov 30 
*+ 16:47:27 CST 2023.

.SUBCKT dffpos Clk D Q 
M_1 Clk_b Clk vdd vdd sky130_fd_pr__pfet_01v8 W='1.26*1u' L=0.15 
+ ad='areap(1.26,sdd)' as='areap(1.26,sdd)' pd='perip(1.26,sdd)' 
+ ps='perip(1.26,sdd)' 
M_2 net_6 net_1 vdd vdd sky130_fd_pr__pfet_01v8 W='0.42*1u' L=0.15 
+ ad='areap(0.42,sdd)' as='areap(0.42,sdd)' pd='perip(0.42,sdd)' 
+ ps='perip(0.42,sdd)' 
M_3 net_4 Clk_b net_6 vdd sky130_fd_pr__pfet_01v8 W='0.42*1u' L=0.15 
+ ad='areap(0.42,sdd)' as='areap(0.42,sdd)' pd='perip(0.42,sdd)' 
+ ps='perip(0.42,sdd)' 
M_4 net_4 Clk net_10 gnd sky130_fd_pr__nfet_01v8 W='0.42*1u' L=0.15 
+ ad='arean(0.42,sdd)' as='arean(0.42,sdd)' pd='perin(0.42,sdd)' 
+ ps='perin(0.42,sdd)' 
M_5 Clk_b Clk gnd gnd sky130_fd_pr__nfet_01v8 W='0.84*1u' L=0.15 
+ ad='arean(0.84,sdd)' as='arean(0.84,sdd)' pd='perin(0.84,sdd)' 
+ ps='perin(0.84,sdd)' 
M_6 net_10 net_1 gnd gnd sky130_fd_pr__nfet_01v8 W='0.42*1u' L=0.15 
+ ad='arean(0.42,sdd)' as='arean(0.42,sdd)' pd='perin(0.42,sdd)' 
+ ps='perin(0.42,sdd)' 
M_7 net_1 net_4 vdd vdd sky130_fd_pr__pfet_01v8 W='0.42*1u' L=0.15 
+ ad='areap(0.42,sdd)' as='areap(0.42,sdd)' pd='perip(0.42,sdd)' 
+ ps='perip(0.42,sdd)' 
M_8 net_1 net_4 gnd gnd sky130_fd_pr__nfet_01v8 W='0.42*1u' L=0.15 
+ ad='arean(0.42,sdd)' as='arean(0.42,sdd)' pd='perin(0.42,sdd)' 
+ ps='perin(0.42,sdd)' 
M_9 net_4 Clk_b net_2 gnd sky130_fd_pr__nfet_01v8 W='0.42*1u' L=0.15 
+ ad='arean(0.42,sdd)' as='arean(0.42,sdd)' pd='perin(0.42,sdd)' 
+ ps='perin(0.42,sdd)' 
M_10 net_2 D gnd gnd sky130_fd_pr__nfet_01v8 W='0.42*1u' L=0.15 
+ ad='arean(0.42,sdd)' as='arean(0.42,sdd)' pd='perin(0.42,sdd)' 
+ ps='perin(0.42,sdd)' 
M_11 net_4 Clk net_8 vdd sky130_fd_pr__pfet_01v8 W='0.42*1u' L=0.15 
+ ad='areap(0.42,sdd)' as='areap(0.42,sdd)' pd='perip(0.42,sdd)' 
+ ps='perip(0.42,sdd)' 
M_12 net_8 D vdd vdd sky130_fd_pr__pfet_01v8 W='0.42*1u' L=0.15 
+ ad='areap(0.42,sdd)' as='areap(0.42,sdd)' pd='perip(0.42,sdd)' 
+ ps='perip(0.42,sdd)' 
M_13 net_3 Clk_b net_9 vdd sky130_fd_pr__pfet_01v8 W='0.42*1u' L=0.15 
+ ad='areap(0.42,sdd)' as='areap(0.42,sdd)' pd='perip(0.42,sdd)' 
+ ps='perip(0.42,sdd)' 
M_14 net_3 Clk net_5 gnd sky130_fd_pr__nfet_01v8 W='0.42*1u' L=0.15 
+ ad='arean(0.42,sdd)' as='arean(0.42,sdd)' pd='perin(0.42,sdd)' 
+ ps='perin(0.42,sdd)' 
M_15 net_5 net_1 gnd gnd sky130_fd_pr__nfet_01v8 W='0.42*1u' L=0.15 
+ ad='arean(0.42,sdd)' as='arean(0.42,sdd)' pd='perin(0.42,sdd)' 
+ ps='perin(0.42,sdd)' 
M_16 net_9 net_1 vdd vdd sky130_fd_pr__pfet_01v8 W='0.42*1u' L=0.15 
+ ad='areap(0.42,sdd)' as='areap(0.42,sdd)' pd='perip(0.42,sdd)' 
+ ps='perip(0.42,sdd)' 
M_17 Q net_3 vdd vdd sky130_fd_pr__pfet_01v8 W='0.84*1u' L=0.15 
+ ad='areap(0.84,sdd)' as='areap(0.84,sdd)' pd='perip(0.84,sdd)' 
+ ps='perip(0.84,sdd)' 
M_18 Q net_3 gnd gnd sky130_fd_pr__nfet_01v8 W='0.42*1u' L=0.15 
+ ad='arean(0.42,sdd)' as='arean(0.42,sdd)' pd='perin(0.42,sdd)' 
+ ps='perin(0.42,sdd)' 
M_19 net_7 Q vdd vdd sky130_fd_pr__pfet_01v8 W='0.42*1u' L=0.15 
+ ad='areap(0.42,sdd)' as='areap(0.42,sdd)' pd='perip(0.42,sdd)' 
+ ps='perip(0.42,sdd)' 
M_20 net_3 Clk net_7 vdd sky130_fd_pr__pfet_01v8 W='0.42*1u' L=0.15 
+ ad='areap(0.42,sdd)' as='areap(0.42,sdd)' pd='perip(0.42,sdd)' 
+ ps='perip(0.42,sdd)' 
M_21 net_3 Clk_b net_11 gnd sky130_fd_pr__nfet_01v8 W='0.42*1u' L=0.15 
+ ad='arean(0.42,sdd)' as='arean(0.42,sdd)' pd='perin(0.42,sdd)' 
+ ps='perin(0.42,sdd)' 
M_22 net_11 Q gnd gnd sky130_fd_pr__nfet_01v8 W='0.42*1u' L=0.15 
+ ad='arean(0.42,sdd)' as='arean(0.42,sdd)' pd='perin(0.42,sdd)' 
+ ps='perin(0.42,sdd)' 
.ENDS	$ dffpos

.SUBCKT inv IN OUT 
Mp0 OUT IN Vdd vdd sky130_fd_pr__pfet_01v8 W='6*1u' L=lp_min 
+ ad='areap(6,sdd)' as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
Mn0 OUT IN Gnd gnd sky130_fd_pr__nfet_01v8 W='3*1u' L=ln_min 
+ ad='arean(3,sdd)' as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
.ENDS	$ inv

.SUBCKT mux21 In_0 In_1 Out Sel Sel_bar 
M_1 Out Sel In_1 gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=ln_min 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
M_2 Out Sel_bar In_1 vdd sky130_fd_pr__pfet_01v8 W='1.26*1u' L=lp_min 
+ ad='areap(1.26,sdd)' as='areap(1.26,sdd)' pd='perip(1.26,sdd)' 
+ ps='perip(1.26,sdd)' 
M_3 Out Sel_bar In_0 gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=ln_min 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
M_4 Out Sel In_0 vdd sky130_fd_pr__pfet_01v8 W='1.26*1u' L=lp_min 
+ ad='areap(1.26,sdd)' as='areap(1.26,sdd)' pd='perip(1.26,sdd)' 
+ ps='perip(1.26,sdd)' 
.ENDS	$ mux21

.SUBCKT FA A B CO Cin S 
M_1 net_5 Cin net_7 vdd sky130_fd_pr__pfet_01v8 W='3*1u' L=0.15u 
+ ad='areap(3,sdd)' as='areap(3,sdd)' pd='perip(3,sdd)' ps='perip(3,sdd)' 
M_2 net_7 B vdd vdd sky130_fd_pr__pfet_01v8 W='3*1u' L=0.15u 
+ ad='areap(3,sdd)' as='areap(3,sdd)' pd='perip(3,sdd)' ps='perip(3,sdd)' 
M_3 net_6 A vdd vdd sky130_fd_pr__pfet_01v8 W='3*1u' L=0.15u 
+ ad='areap(3,sdd)' as='areap(3,sdd)' pd='perip(3,sdd)' ps='perip(3,sdd)' 
M_4 net_5 B net_6 vdd sky130_fd_pr__pfet_01v8 W='3*1u' L=0.15u 
+ ad='areap(3,sdd)' as='areap(3,sdd)' pd='perip(3,sdd)' ps='perip(3,sdd)' 
M_5 net_11 A vdd vdd sky130_fd_pr__pfet_01v8 W='3.0*1u' L=0.15u 
+ ad='areap(3.0,sdd)' as='areap(3.0,sdd)' pd='perip(3.0,sdd)' 
+ ps='perip(3.0,sdd)' 
M_6 net_11 B vdd vdd sky130_fd_pr__pfet_01v8 W='3.0*1u' L=0.15u 
+ ad='areap(3.0,sdd)' as='areap(3.0,sdd)' pd='perip(3.0,sdd)' 
+ ps='perip(3.0,sdd)' 
M_7 net_11 Cin vdd vdd sky130_fd_pr__pfet_01v8 W='3.0*1u' L=0.15u 
+ ad='areap(3.0,sdd)' as='areap(3.0,sdd)' pd='perip(3.0,sdd)' 
+ ps='perip(3.0,sdd)' 
M_8 net_10 Cin net_1 vdd sky130_fd_pr__pfet_01v8 W='3.0*1u' L=0.15u 
+ ad='areap(3.0,sdd)' as='areap(3.0,sdd)' pd='perip(3.0,sdd)' 
+ ps='perip(3.0,sdd)' 
M_9 net_1 B net_2 vdd sky130_fd_pr__pfet_01v8 W='3.0*1u' L=0.15u 
+ ad='areap(3.0,sdd)' as='areap(3.0,sdd)' pd='perip(3.0,sdd)' 
+ ps='perip(3.0,sdd)' 
M_10 net_2 A vdd vdd sky130_fd_pr__pfet_01v8 W='3.0*1u' L=0.15u 
+ ad='areap(3.0,sdd)' as='areap(3.0,sdd)' pd='perip(3.0,sdd)' 
+ ps='perip(3.0,sdd)' 
M_11 net_10 net_5 net_11 vdd sky130_fd_pr__pfet_01v8 W='3.0*1u' L=0.15u 
+ ad='areap(3.0,sdd)' as='areap(3.0,sdd)' pd='perip(3.0,sdd)' 
+ ps='perip(3.0,sdd)' 
M_12 net_7 A vdd vdd sky130_fd_pr__pfet_01v8 W='3.0*1u' L=0.15u 
+ ad='areap(3.0,sdd)' as='areap(3.0,sdd)' pd='perip(3.0,sdd)' 
+ ps='perip(3.0,sdd)' 
M_13 net_5 Cin net_3 gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=0.15u 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
M_14 net_3 A gnd gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=0.15u 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
M_15 net_3 B gnd gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=0.15u 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
M_16 net_4 A gnd gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=0.15u 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
M_17 net_5 B net_4 gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=0.15u 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
M_18 net_9 A gnd gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=0.15u 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
M_19 net_9 B gnd gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=0.15u 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
M_20 net_9 Cin gnd gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=0.15u 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
M_21 net_10 net_5 net_9 gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=0.15u 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
M_22 net_10 Cin net_12 gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=0.15u 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
M_23 net_12 B net_8 gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=0.15u 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
M_24 net_8 A gnd gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=0.15u 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
M_25 CO net_5 vdd vdd sky130_fd_pr__pfet_01v8 W='3*1u' L=0.15u 
+ ad='areap(3,sdd)' as='areap(3,sdd)' pd='perip(3,sdd)' ps='perip(3,sdd)' 
M_26 CO net_5 gnd gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=0.15u 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
M_27 S net_10 vdd vdd sky130_fd_pr__pfet_01v8 W='3*1u' L=0.15u 
+ ad='areap(3,sdd)' as='areap(3,sdd)' pd='perip(3,sdd)' ps='perip(3,sdd)' 
M_28 S net_10 gnd gnd sky130_fd_pr__nfet_01v8 W='0.52*1u' L=0.15u 
+ ad='arean(0.52,sdd)' as='arean(0.52,sdd)' pd='perin(0.52,sdd)' 
+ ps='perin(0.52,sdd)' 
.ENDS	$ FA

.SUBCKT bit1a A B Cin Cout EN Out clk 
Xdffpos clk net_3 Out dffpos 
Xinv EN net_2 inv 
Xmux21 Out net_1 net_3 EN net_2 mux21 
XFA A B Cout Cin net_1 FA 
.ENDS	$ bit1a

* start main CELL top
* .SUBCKT top A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] B[0] B[1] B[2] 
*+ B[3] B[4] B[5] B[6] B[7] Z[0] Z[1] Z[2] Z[3] Z[4] Z[5] Z[6] Z[7] cin 
*+ clk en 
Xbit1a A[0] B[0] cin c[1] en Z[0] clk bit1a 
Xbit1a_1 A[1] B[1] c[1] c[2] en Z[1] clk bit1a 
Xbit1a_2 A[2] B[2] c[2] c[3] en Z[2] clk bit1a 
Xbit1a_3 A[3] B[3] c[3] c[4] en Z[3] clk bit1a 
Xbit1a_4 A[7] B[7] c[7] Z[8] en Z[7] clk bit1a 
Xbit1a_5 A[6] B[6] c[6] c[7] en Z[6] clk bit1a 
Xbit1a_6 A[5] B[5] c[5] c[6] en Z[5] clk bit1a 
Xbit1a_7 A[4] B[4] c[4] c[5] en Z[4] clk bit1a 
* .ENDS	$ top

.GLOBAL gnd vdd

.END


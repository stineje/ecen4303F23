magic
tech scmos
timestamp 1084294368
<< nwell >>
rect 20 740 280 1000
rect 15 604 286 652
rect 14 475 286 604
rect 14 425 285 475
rect 142 424 285 425
rect -6 253 303 338
rect -3 249 303 253
rect -3 11 11 249
rect 286 11 303 249
rect -3 -3 303 11
<< pwell >>
rect -3 654 303 673
rect -3 423 14 654
rect 114 423 186 424
rect 286 423 303 654
rect -3 407 303 423
rect -3 389 9 407
rect 290 389 303 407
rect -3 351 162 389
rect 186 351 303 389
rect -3 338 303 351
rect 11 11 284 249
<< ntransistor >>
rect 19 353 21 383
rect 27 353 29 383
rect 44 353 46 383
rect 52 353 54 383
rect 60 353 62 383
rect 68 353 70 383
rect 76 353 78 383
rect 84 353 86 383
rect 92 353 94 383
rect 100 353 102 383
rect 108 353 110 383
rect 116 353 118 383
rect 124 353 126 383
rect 132 353 134 383
rect 140 353 142 383
rect 148 353 150 383
rect 198 353 200 383
rect 206 353 208 383
rect 214 353 216 383
rect 222 353 224 383
rect 230 353 232 383
rect 238 353 240 383
rect 246 353 248 383
rect 254 353 256 383
rect 262 353 264 383
rect 270 353 272 383
rect 278 353 280 383
rect 286 353 288 383
rect 38 216 138 219
rect 38 171 138 174
rect 38 150 138 153
rect 38 106 138 109
rect 38 85 138 88
rect 38 41 138 44
rect 162 216 262 219
rect 162 171 262 174
rect 162 150 262 153
rect 162 106 262 109
rect 162 85 262 88
rect 162 41 262 44
<< ptransistor >>
rect 38 624 138 627
rect 38 580 138 583
rect 38 559 138 562
rect 38 516 138 519
rect 38 495 138 498
rect 38 451 138 454
rect 162 624 262 627
rect 162 580 262 583
rect 162 559 262 562
rect 162 516 262 519
rect 162 495 262 498
rect 162 451 262 454
rect 19 269 21 321
rect 27 269 29 321
rect 44 269 46 321
rect 52 269 54 321
rect 60 269 62 321
rect 68 269 70 321
rect 76 269 78 321
rect 84 269 86 321
rect 92 269 94 321
rect 100 269 102 321
rect 108 269 110 321
rect 116 269 118 321
rect 124 269 126 321
rect 132 269 134 321
rect 140 269 142 321
rect 148 269 150 321
rect 198 269 200 321
rect 206 269 208 321
rect 214 269 216 321
rect 222 269 224 321
rect 230 269 232 321
rect 238 269 240 321
rect 246 269 248 321
rect 254 269 256 321
rect 262 269 264 321
rect 270 269 272 321
rect 278 269 280 321
rect 286 269 288 321
<< ndiffusion >>
rect 13 380 19 383
rect 13 361 14 380
rect 18 361 19 380
rect 13 353 19 361
rect 21 380 27 383
rect 21 376 22 380
rect 26 376 27 380
rect 21 370 27 376
rect 21 366 22 370
rect 26 366 27 370
rect 21 360 27 366
rect 21 356 22 360
rect 26 356 27 360
rect 21 353 27 356
rect 29 379 35 383
rect 29 355 30 379
rect 34 355 35 379
rect 29 353 35 355
rect 38 379 44 383
rect 38 360 39 379
rect 43 360 44 379
rect 38 353 44 360
rect 46 378 52 383
rect 46 374 47 378
rect 51 374 52 378
rect 46 368 52 374
rect 46 364 47 368
rect 51 364 52 368
rect 46 358 52 364
rect 46 354 47 358
rect 51 354 52 358
rect 46 353 52 354
rect 54 379 60 383
rect 54 355 55 379
rect 59 355 60 379
rect 54 353 60 355
rect 62 378 68 383
rect 62 374 63 378
rect 67 374 68 378
rect 62 368 68 374
rect 62 364 63 368
rect 67 364 68 368
rect 62 358 68 364
rect 62 354 63 358
rect 67 354 68 358
rect 62 353 68 354
rect 70 379 76 383
rect 70 355 71 379
rect 75 355 76 379
rect 70 353 76 355
rect 78 378 84 383
rect 78 374 79 378
rect 83 374 84 378
rect 78 368 84 374
rect 78 364 79 368
rect 83 364 84 368
rect 78 358 84 364
rect 78 354 79 358
rect 83 354 84 358
rect 78 353 84 354
rect 86 379 92 383
rect 86 355 87 379
rect 91 355 92 379
rect 86 353 92 355
rect 94 378 100 383
rect 94 374 95 378
rect 99 374 100 378
rect 94 368 100 374
rect 94 364 95 368
rect 99 364 100 368
rect 94 358 100 364
rect 94 354 95 358
rect 99 354 100 358
rect 94 353 100 354
rect 102 380 108 383
rect 102 356 103 380
rect 107 356 108 380
rect 102 353 108 356
rect 110 378 116 383
rect 110 374 111 378
rect 115 374 116 378
rect 110 368 116 374
rect 110 364 111 368
rect 115 364 116 368
rect 110 358 116 364
rect 110 354 111 358
rect 115 354 116 358
rect 110 353 116 354
rect 118 379 124 383
rect 118 365 119 379
rect 123 365 124 379
rect 118 353 124 365
rect 126 378 132 383
rect 126 354 127 378
rect 131 354 132 378
rect 126 353 132 354
rect 134 379 140 383
rect 134 365 135 379
rect 139 365 140 379
rect 134 359 140 365
rect 134 355 135 359
rect 139 355 140 359
rect 134 353 140 355
rect 142 379 148 383
rect 142 360 143 379
rect 147 360 148 379
rect 142 353 148 360
rect 150 382 156 383
rect 150 353 151 382
rect 155 353 156 382
rect 192 380 198 383
rect 192 376 193 380
rect 197 376 198 380
rect 192 370 198 376
rect 192 366 193 370
rect 197 366 198 370
rect 192 360 198 366
rect 192 356 193 360
rect 197 356 198 360
rect 192 353 198 356
rect 200 380 206 383
rect 200 356 201 380
rect 205 356 206 380
rect 200 353 206 356
rect 208 374 214 383
rect 208 365 209 374
rect 213 365 214 374
rect 208 358 214 365
rect 208 354 209 358
rect 213 354 214 358
rect 208 353 214 354
rect 216 380 222 383
rect 216 356 217 380
rect 221 356 222 380
rect 216 353 222 356
rect 224 380 230 383
rect 224 376 225 380
rect 229 376 230 380
rect 224 370 230 376
rect 224 366 225 370
rect 229 366 230 370
rect 224 360 230 366
rect 224 356 225 360
rect 229 356 230 360
rect 224 353 230 356
rect 232 380 238 383
rect 232 356 233 380
rect 237 356 238 380
rect 232 353 238 356
rect 240 380 246 383
rect 240 376 241 380
rect 245 376 246 380
rect 240 370 246 376
rect 240 366 241 370
rect 245 366 246 370
rect 240 360 246 366
rect 240 356 241 360
rect 245 356 246 360
rect 240 353 246 356
rect 248 380 254 383
rect 248 356 249 380
rect 253 356 254 380
rect 248 353 254 356
rect 256 380 262 383
rect 256 376 257 380
rect 261 376 262 380
rect 256 370 262 376
rect 256 366 257 370
rect 261 366 262 370
rect 256 360 262 366
rect 256 356 257 360
rect 261 356 262 360
rect 256 353 262 356
rect 264 380 270 383
rect 264 356 265 380
rect 269 356 270 380
rect 264 353 270 356
rect 272 380 278 383
rect 272 376 273 380
rect 277 376 278 380
rect 272 370 278 376
rect 272 366 273 370
rect 277 366 278 370
rect 272 360 278 366
rect 272 356 273 360
rect 277 356 278 360
rect 272 353 278 356
rect 280 380 286 383
rect 280 356 281 380
rect 285 356 286 380
rect 280 353 286 356
rect 288 380 293 383
rect 288 376 289 380
rect 288 370 293 376
rect 288 366 289 370
rect 288 360 293 366
rect 288 356 289 360
rect 288 353 293 356
rect 47 350 50 353
rect 63 350 67 353
rect 79 350 83 353
rect 111 350 115 353
rect 192 350 197 353
rect 209 350 213 353
rect 225 350 228 353
rect 241 350 245 353
rect 257 350 261 353
rect 273 350 276 353
rect 289 350 293 353
rect 38 227 138 228
rect 38 223 54 227
rect 63 223 69 227
rect 78 223 84 227
rect 93 223 99 227
rect 108 223 114 227
rect 118 223 138 227
rect 38 219 138 223
rect 38 200 138 216
rect 38 196 56 200
rect 120 196 138 200
rect 38 194 138 196
rect 38 190 56 194
rect 120 190 138 194
rect 38 174 138 190
rect 38 167 138 171
rect 38 163 55 167
rect 64 163 70 167
rect 79 163 85 167
rect 94 163 100 167
rect 109 163 115 167
rect 119 163 138 167
rect 38 161 138 163
rect 38 157 55 161
rect 64 157 70 161
rect 79 157 85 161
rect 94 157 100 161
rect 109 157 115 161
rect 119 157 138 161
rect 38 153 138 157
rect 38 134 138 150
rect 38 125 56 134
rect 120 125 138 134
rect 38 109 138 125
rect 38 102 138 106
rect 38 98 54 102
rect 63 98 69 102
rect 78 98 84 102
rect 93 98 99 102
rect 108 98 114 102
rect 118 98 138 102
rect 38 96 138 98
rect 38 92 54 96
rect 63 92 69 96
rect 78 92 84 96
rect 93 92 99 96
rect 108 92 114 96
rect 118 92 138 96
rect 38 88 138 92
rect 38 69 138 85
rect 38 60 56 69
rect 120 60 138 69
rect 38 44 138 60
rect 162 227 262 228
rect 162 223 182 227
rect 191 223 197 227
rect 206 223 212 227
rect 221 223 227 227
rect 236 223 242 227
rect 246 223 262 227
rect 162 219 262 223
rect 38 37 138 41
rect 38 33 39 37
rect 43 33 53 37
rect 57 33 59 37
rect 118 33 138 37
rect 38 32 138 33
rect 38 31 43 32
rect 162 200 262 216
rect 162 196 180 200
rect 244 196 262 200
rect 162 194 262 196
rect 162 190 180 194
rect 244 190 262 194
rect 162 174 262 190
rect 162 167 262 171
rect 162 163 181 167
rect 190 163 196 167
rect 205 163 211 167
rect 220 163 226 167
rect 235 163 241 167
rect 245 163 262 167
rect 162 161 262 163
rect 162 157 181 161
rect 190 157 196 161
rect 205 157 211 161
rect 220 157 226 161
rect 235 157 241 161
rect 245 157 262 161
rect 162 153 262 157
rect 162 134 262 150
rect 162 125 180 134
rect 244 125 262 134
rect 162 109 262 125
rect 162 102 262 106
rect 162 98 182 102
rect 191 98 197 102
rect 206 98 212 102
rect 221 98 227 102
rect 236 98 242 102
rect 246 98 262 102
rect 162 96 262 98
rect 162 92 182 96
rect 191 92 197 96
rect 206 92 212 96
rect 221 92 227 96
rect 236 92 242 96
rect 246 92 262 96
rect 162 88 262 92
rect 162 69 262 85
rect 162 60 180 69
rect 244 60 262 69
rect 162 44 262 60
rect 162 37 262 41
rect 162 33 182 37
rect 246 33 262 37
rect 162 32 262 33
<< pdiffusion >>
rect 36 634 140 636
rect 36 630 45 634
rect 54 630 56 634
rect 60 630 66 634
rect 75 630 81 634
rect 90 630 96 634
rect 105 630 111 634
rect 115 630 140 634
rect 38 629 141 630
rect 38 627 138 629
rect 38 608 138 624
rect 38 599 56 608
rect 120 599 138 608
rect 38 583 138 599
rect 38 576 138 580
rect 38 572 61 576
rect 70 572 76 576
rect 85 572 91 576
rect 100 572 106 576
rect 115 572 138 576
rect 38 570 138 572
rect 38 566 61 570
rect 70 566 76 570
rect 85 566 91 570
rect 100 566 106 570
rect 115 566 138 570
rect 38 562 138 566
rect 38 543 138 559
rect 38 534 56 543
rect 120 534 138 543
rect 38 519 138 534
rect 38 512 138 516
rect 38 508 61 512
rect 70 508 76 512
rect 85 508 91 512
rect 100 508 106 512
rect 115 508 138 512
rect 38 506 138 508
rect 38 502 61 506
rect 70 502 76 506
rect 85 502 91 506
rect 100 502 106 506
rect 115 502 138 506
rect 38 498 138 502
rect 38 479 138 495
rect 38 470 56 479
rect 120 470 138 479
rect 38 454 138 470
rect 160 634 264 636
rect 160 630 183 634
rect 187 630 193 634
rect 202 630 208 634
rect 217 630 223 634
rect 232 630 238 634
rect 242 630 244 634
rect 253 630 264 634
rect 159 629 262 630
rect 162 627 262 629
rect 38 447 138 451
rect 38 443 61 447
rect 70 443 76 447
rect 85 443 91 447
rect 100 443 106 447
rect 115 443 138 447
rect 38 442 138 443
rect 162 608 262 624
rect 162 599 180 608
rect 244 599 262 608
rect 162 583 262 599
rect 162 576 262 580
rect 162 572 184 576
rect 193 572 199 576
rect 208 572 214 576
rect 223 572 229 576
rect 238 572 262 576
rect 162 570 262 572
rect 162 566 184 570
rect 193 566 199 570
rect 208 566 214 570
rect 223 566 229 570
rect 238 566 262 570
rect 162 562 262 566
rect 162 543 262 559
rect 162 534 180 543
rect 244 534 262 543
rect 162 519 262 534
rect 162 512 262 516
rect 162 508 183 512
rect 192 508 198 512
rect 207 508 213 512
rect 222 508 228 512
rect 237 508 262 512
rect 162 506 262 508
rect 162 502 183 506
rect 192 502 198 506
rect 207 502 213 506
rect 222 502 228 506
rect 237 502 262 506
rect 162 498 262 502
rect 162 479 262 495
rect 162 470 180 479
rect 244 470 262 479
rect 162 454 262 470
rect 162 447 262 451
rect 162 443 184 447
rect 193 443 199 447
rect 208 443 214 447
rect 223 443 229 447
rect 238 443 262 447
rect 162 442 262 443
rect 63 321 67 324
rect 79 321 83 324
rect 111 321 115 324
rect 192 321 197 324
rect 209 321 213 324
rect 225 321 228 324
rect 241 321 245 324
rect 257 321 261 324
rect 273 321 276 324
rect 289 321 293 324
rect 13 314 19 321
rect 13 270 14 314
rect 18 270 19 314
rect 13 269 19 270
rect 21 320 27 321
rect 21 316 22 320
rect 26 316 27 320
rect 21 310 27 316
rect 21 306 22 310
rect 26 306 27 310
rect 21 300 27 306
rect 21 296 22 300
rect 26 296 27 300
rect 21 290 27 296
rect 21 286 22 290
rect 26 286 27 290
rect 21 280 27 286
rect 21 276 22 280
rect 26 276 27 280
rect 21 269 27 276
rect 29 319 35 321
rect 29 270 30 319
rect 34 270 35 319
rect 29 269 35 270
rect 38 314 44 321
rect 38 270 39 314
rect 43 270 44 314
rect 38 269 44 270
rect 46 320 52 321
rect 46 316 47 320
rect 51 316 52 320
rect 46 310 52 316
rect 46 306 47 310
rect 51 306 52 310
rect 46 300 52 306
rect 46 296 47 300
rect 51 296 52 300
rect 46 290 52 296
rect 46 286 47 290
rect 51 286 52 290
rect 46 280 52 286
rect 46 276 47 280
rect 51 276 52 280
rect 46 269 52 276
rect 54 319 60 321
rect 54 270 55 319
rect 59 270 60 319
rect 54 269 60 270
rect 62 316 68 321
rect 62 312 63 316
rect 67 312 68 316
rect 62 306 68 312
rect 62 302 63 306
rect 67 302 68 306
rect 62 296 68 302
rect 62 292 63 296
rect 67 292 68 296
rect 62 286 68 292
rect 62 282 63 286
rect 67 282 68 286
rect 62 276 68 282
rect 62 272 63 276
rect 67 272 68 276
rect 62 269 68 272
rect 70 319 76 321
rect 70 270 71 319
rect 75 270 76 319
rect 70 269 76 270
rect 78 316 84 321
rect 78 312 79 316
rect 83 312 84 316
rect 78 306 84 312
rect 78 302 79 306
rect 83 302 84 306
rect 78 296 84 302
rect 78 292 79 296
rect 83 292 84 296
rect 78 286 84 292
rect 78 282 79 286
rect 83 282 84 286
rect 78 276 84 282
rect 78 272 79 276
rect 83 272 84 276
rect 78 269 84 272
rect 86 320 92 321
rect 86 271 87 320
rect 91 271 92 320
rect 86 269 92 271
rect 94 316 100 321
rect 94 312 95 316
rect 99 312 100 316
rect 94 306 100 312
rect 94 302 95 306
rect 99 302 100 306
rect 94 296 100 302
rect 94 292 95 296
rect 99 292 100 296
rect 94 286 100 292
rect 94 282 95 286
rect 99 282 100 286
rect 94 276 100 282
rect 94 272 95 276
rect 99 272 100 276
rect 94 269 100 272
rect 102 319 108 321
rect 102 270 103 319
rect 107 270 108 319
rect 102 269 108 270
rect 110 320 116 321
rect 110 316 111 320
rect 115 316 116 320
rect 110 310 116 316
rect 110 306 111 310
rect 115 306 116 310
rect 110 300 116 306
rect 110 296 111 300
rect 115 296 116 300
rect 110 290 116 296
rect 110 286 111 290
rect 115 286 116 290
rect 110 280 116 286
rect 110 276 111 280
rect 115 276 116 280
rect 110 269 116 276
rect 118 320 124 321
rect 118 271 119 320
rect 123 271 124 320
rect 118 269 124 271
rect 126 311 132 321
rect 126 272 127 311
rect 131 272 132 311
rect 126 269 132 272
rect 134 320 140 321
rect 134 316 135 320
rect 139 316 140 320
rect 134 307 140 316
rect 134 278 135 307
rect 139 278 140 307
rect 134 269 140 278
rect 142 320 148 321
rect 142 271 143 320
rect 147 271 148 320
rect 142 269 148 271
rect 150 309 156 321
rect 150 270 151 309
rect 155 270 156 309
rect 150 269 156 270
rect 192 316 198 321
rect 192 312 193 316
rect 197 312 198 316
rect 192 306 198 312
rect 192 302 193 306
rect 197 302 198 306
rect 192 291 198 302
rect 192 282 193 291
rect 197 282 198 291
rect 192 276 198 282
rect 192 272 193 276
rect 197 272 198 276
rect 192 269 198 272
rect 200 316 206 321
rect 200 272 201 316
rect 205 272 206 316
rect 200 269 206 272
rect 208 316 214 321
rect 208 312 209 316
rect 213 312 214 316
rect 208 306 214 312
rect 208 302 209 306
rect 213 302 214 306
rect 208 291 214 302
rect 208 282 209 291
rect 213 282 214 291
rect 208 276 214 282
rect 208 272 209 276
rect 213 272 214 276
rect 208 269 214 272
rect 216 316 222 321
rect 216 272 217 316
rect 221 272 222 316
rect 216 269 222 272
rect 224 316 230 321
rect 224 312 225 316
rect 229 312 230 316
rect 224 306 230 312
rect 224 302 225 306
rect 229 302 230 306
rect 224 291 230 302
rect 224 282 225 291
rect 229 282 230 291
rect 224 276 230 282
rect 224 272 225 276
rect 229 272 230 276
rect 224 269 230 272
rect 232 316 238 321
rect 232 272 233 316
rect 237 272 238 316
rect 232 269 238 272
rect 240 316 246 321
rect 240 312 241 316
rect 245 312 246 316
rect 240 306 246 312
rect 240 302 241 306
rect 245 302 246 306
rect 240 291 246 302
rect 240 282 241 291
rect 245 282 246 291
rect 240 276 246 282
rect 240 272 241 276
rect 245 272 246 276
rect 240 269 246 272
rect 248 316 254 321
rect 248 272 249 316
rect 253 272 254 316
rect 248 269 254 272
rect 256 316 262 321
rect 256 312 257 316
rect 261 312 262 316
rect 256 306 262 312
rect 256 302 257 306
rect 261 302 262 306
rect 256 291 262 302
rect 256 282 257 291
rect 261 282 262 291
rect 256 276 262 282
rect 256 272 257 276
rect 261 272 262 276
rect 256 269 262 272
rect 264 316 270 321
rect 264 272 265 316
rect 269 272 270 316
rect 264 269 270 272
rect 272 316 278 321
rect 272 312 273 316
rect 277 312 278 316
rect 272 306 278 312
rect 272 302 273 306
rect 277 302 278 306
rect 272 291 278 302
rect 272 282 273 291
rect 277 282 278 291
rect 272 276 278 282
rect 272 272 273 276
rect 277 272 278 276
rect 272 269 278 272
rect 280 316 286 321
rect 280 272 281 316
rect 285 272 286 316
rect 280 269 286 272
rect 288 316 293 321
rect 288 269 289 316
rect 79 266 83 269
rect 192 266 197 269
rect 241 266 245 269
<< ndcontact >>
rect 14 361 18 380
rect 22 376 26 380
rect 22 366 26 370
rect 22 356 26 360
rect 30 355 34 379
rect 39 360 43 379
rect 47 374 51 378
rect 47 364 51 368
rect 47 354 51 358
rect 55 355 59 379
rect 63 374 67 378
rect 63 364 67 368
rect 63 354 67 358
rect 71 355 75 379
rect 79 374 83 378
rect 79 364 83 368
rect 79 354 83 358
rect 87 355 91 379
rect 95 374 99 378
rect 95 364 99 368
rect 95 354 99 358
rect 103 356 107 380
rect 111 374 115 378
rect 111 364 115 368
rect 111 354 115 358
rect 119 365 123 379
rect 127 354 131 378
rect 135 365 139 379
rect 135 355 139 359
rect 143 360 147 379
rect 151 353 155 382
rect 193 376 197 380
rect 193 366 197 370
rect 193 356 197 360
rect 201 356 205 380
rect 209 365 213 374
rect 209 354 213 358
rect 217 356 221 380
rect 225 376 229 380
rect 225 366 229 370
rect 225 356 229 360
rect 233 356 237 380
rect 241 376 245 380
rect 241 366 245 370
rect 241 356 245 360
rect 249 356 253 380
rect 257 376 261 380
rect 257 366 261 370
rect 257 356 261 360
rect 265 356 269 380
rect 273 376 277 380
rect 273 366 277 370
rect 273 356 277 360
rect 281 356 285 380
rect 289 376 293 380
rect 289 366 293 370
rect 289 356 293 360
rect 54 223 63 227
rect 69 223 78 227
rect 84 223 93 227
rect 99 223 108 227
rect 114 223 118 227
rect 56 196 120 200
rect 56 190 120 194
rect 55 163 64 167
rect 70 163 79 167
rect 85 163 94 167
rect 100 163 109 167
rect 115 163 119 167
rect 55 157 64 161
rect 70 157 79 161
rect 85 157 94 161
rect 100 157 109 161
rect 115 157 119 161
rect 56 125 120 134
rect 54 98 63 102
rect 69 98 78 102
rect 84 98 93 102
rect 99 98 108 102
rect 114 98 118 102
rect 54 92 63 96
rect 69 92 78 96
rect 84 92 93 96
rect 99 92 108 96
rect 114 92 118 96
rect 56 60 120 69
rect 182 223 191 227
rect 197 223 206 227
rect 212 223 221 227
rect 227 223 236 227
rect 242 223 246 227
rect 39 33 43 37
rect 53 33 57 37
rect 59 33 118 37
rect 180 196 244 200
rect 180 190 244 194
rect 181 163 190 167
rect 196 163 205 167
rect 211 163 220 167
rect 226 163 235 167
rect 241 163 245 167
rect 181 157 190 161
rect 196 157 205 161
rect 211 157 220 161
rect 226 157 235 161
rect 241 157 245 161
rect 180 125 244 134
rect 182 98 191 102
rect 197 98 206 102
rect 212 98 221 102
rect 227 98 236 102
rect 242 98 246 102
rect 182 92 191 96
rect 197 92 206 96
rect 212 92 221 96
rect 227 92 236 96
rect 242 92 246 96
rect 180 60 244 69
rect 182 33 246 37
<< pdcontact >>
rect 45 630 54 634
rect 56 630 60 634
rect 66 630 75 634
rect 81 630 90 634
rect 96 630 105 634
rect 111 630 115 634
rect 56 599 120 608
rect 61 572 70 576
rect 76 572 85 576
rect 91 572 100 576
rect 106 572 115 576
rect 61 566 70 570
rect 76 566 85 570
rect 91 566 100 570
rect 106 566 115 570
rect 56 534 120 543
rect 61 508 70 512
rect 76 508 85 512
rect 91 508 100 512
rect 106 508 115 512
rect 61 502 70 506
rect 76 502 85 506
rect 91 502 100 506
rect 106 502 115 506
rect 56 470 120 479
rect 183 630 187 634
rect 193 630 202 634
rect 208 630 217 634
rect 223 630 232 634
rect 238 630 242 634
rect 244 630 253 634
rect 61 443 70 447
rect 76 443 85 447
rect 91 443 100 447
rect 106 443 115 447
rect 180 599 244 608
rect 184 572 193 576
rect 199 572 208 576
rect 214 572 223 576
rect 229 572 238 576
rect 184 566 193 570
rect 199 566 208 570
rect 214 566 223 570
rect 229 566 238 570
rect 180 534 244 543
rect 183 508 192 512
rect 198 508 207 512
rect 213 508 222 512
rect 228 508 237 512
rect 183 502 192 506
rect 198 502 207 506
rect 213 502 222 506
rect 228 502 237 506
rect 180 470 244 479
rect 184 443 193 447
rect 199 443 208 447
rect 214 443 223 447
rect 229 443 238 447
rect 14 270 18 314
rect 22 316 26 320
rect 22 306 26 310
rect 22 296 26 300
rect 22 286 26 290
rect 22 276 26 280
rect 30 270 34 319
rect 39 270 43 314
rect 47 316 51 320
rect 47 306 51 310
rect 47 296 51 300
rect 47 286 51 290
rect 47 276 51 280
rect 55 270 59 319
rect 63 312 67 316
rect 63 302 67 306
rect 63 292 67 296
rect 63 282 67 286
rect 63 272 67 276
rect 71 270 75 319
rect 79 312 83 316
rect 79 302 83 306
rect 79 292 83 296
rect 79 282 83 286
rect 79 272 83 276
rect 87 271 91 320
rect 95 312 99 316
rect 95 302 99 306
rect 95 292 99 296
rect 95 282 99 286
rect 95 272 99 276
rect 103 270 107 319
rect 111 316 115 320
rect 111 306 115 310
rect 111 296 115 300
rect 111 286 115 290
rect 111 276 115 280
rect 119 271 123 320
rect 127 272 131 311
rect 135 316 139 320
rect 135 278 139 307
rect 143 271 147 320
rect 151 270 155 309
rect 193 312 197 316
rect 193 302 197 306
rect 193 282 197 291
rect 193 272 197 276
rect 201 272 205 316
rect 209 312 213 316
rect 209 302 213 306
rect 209 282 213 291
rect 209 272 213 276
rect 217 272 221 316
rect 225 312 229 316
rect 225 302 229 306
rect 225 282 229 291
rect 225 272 229 276
rect 233 272 237 316
rect 241 312 245 316
rect 241 302 245 306
rect 241 282 245 291
rect 241 272 245 276
rect 249 272 253 316
rect 257 312 261 316
rect 257 302 261 306
rect 257 282 261 291
rect 257 272 261 276
rect 265 272 269 316
rect 273 312 277 316
rect 273 302 277 306
rect 273 282 277 291
rect 273 272 277 276
rect 281 272 285 316
rect 289 257 293 316
<< psubstratepdiff >>
rect 0 667 300 670
rect 0 658 1 667
rect 115 658 184 667
rect 298 658 300 667
rect 0 657 300 658
rect 0 654 11 657
rect 0 415 1 654
rect 10 420 11 654
rect 289 656 300 657
rect 117 420 147 421
rect 153 420 183 421
rect 289 420 290 656
rect 10 419 290 420
rect 10 415 15 419
rect 0 410 15 415
rect 29 410 39 419
rect 113 410 148 419
rect 152 410 184 419
rect 288 412 290 419
rect 299 412 300 656
rect 288 410 300 412
rect 0 407 6 410
rect 0 343 1 407
rect 5 348 6 407
rect 293 406 300 410
rect 293 402 295 406
rect 299 402 300 406
rect 293 396 300 402
rect 293 392 295 396
rect 299 392 300 396
rect 293 386 300 392
rect 293 382 295 386
rect 299 382 300 386
rect 293 376 300 382
rect 293 372 295 376
rect 299 372 300 376
rect 293 366 300 372
rect 293 362 295 366
rect 299 362 300 366
rect 293 356 300 362
rect 5 345 7 348
rect 15 347 23 348
rect 15 345 17 347
rect 5 343 17 345
rect 21 345 23 347
rect 47 347 50 350
rect 31 346 50 347
rect 31 345 38 346
rect 21 343 38 345
rect 0 342 38 343
rect 42 342 45 346
rect 49 344 50 346
rect 63 347 67 350
rect 79 347 83 350
rect 111 348 115 350
rect 63 346 84 347
rect 97 347 135 348
rect 63 344 64 346
rect 49 342 64 344
rect 83 345 84 346
rect 97 345 99 347
rect 83 343 99 345
rect 103 343 108 347
rect 112 343 124 347
rect 128 345 135 347
rect 192 348 197 350
rect 209 348 213 350
rect 225 348 228 350
rect 148 347 228 348
rect 148 346 223 347
rect 148 345 194 346
rect 128 343 194 345
rect 83 342 194 343
rect 213 343 223 346
rect 227 345 228 347
rect 241 348 245 350
rect 257 348 261 350
rect 273 348 276 350
rect 241 346 276 348
rect 293 352 295 356
rect 299 352 300 356
rect 293 350 300 352
rect 289 346 300 350
rect 241 345 242 346
rect 227 343 242 345
rect 213 342 242 343
rect 251 342 257 346
rect 261 342 271 346
rect 275 345 276 346
rect 289 345 290 346
rect 275 342 290 345
rect 299 342 300 346
rect 0 341 300 342
rect 14 243 281 246
rect 14 241 270 243
rect 14 240 53 241
rect 14 236 17 240
rect 36 237 53 240
rect 117 239 182 241
rect 117 237 148 239
rect 36 236 148 237
rect 14 233 148 236
rect 14 232 54 233
rect 14 228 17 232
rect 26 230 54 232
rect 26 228 30 230
rect 14 222 30 228
rect 14 208 17 222
rect 26 208 30 222
rect 38 229 54 230
rect 63 229 69 233
rect 78 229 84 233
rect 93 229 99 233
rect 108 229 114 233
rect 118 230 148 233
rect 152 237 182 239
rect 246 237 270 241
rect 152 233 270 237
rect 152 230 182 233
rect 118 229 138 230
rect 38 228 138 229
rect 143 224 157 230
rect 14 202 30 208
rect 14 188 17 202
rect 26 188 30 202
rect 14 182 30 188
rect 14 168 17 182
rect 26 168 30 182
rect 14 162 30 168
rect 14 148 17 162
rect 26 148 30 162
rect 14 142 30 148
rect 14 128 17 142
rect 26 128 30 142
rect 14 122 30 128
rect 14 108 17 122
rect 26 108 30 122
rect 14 102 30 108
rect 14 88 17 102
rect 26 88 30 102
rect 14 82 30 88
rect 14 68 17 82
rect 26 68 30 82
rect 14 62 30 68
rect 14 48 17 62
rect 26 48 30 62
rect 14 42 30 48
rect 14 33 17 42
rect 26 33 30 42
rect 143 215 148 224
rect 152 215 157 224
rect 162 229 182 230
rect 191 229 197 233
rect 206 229 212 233
rect 221 229 227 233
rect 236 229 242 233
rect 246 230 270 233
rect 246 229 262 230
rect 162 228 262 229
rect 274 229 276 243
rect 143 209 157 215
rect 143 200 148 209
rect 152 200 157 209
rect 143 194 157 200
rect 143 185 148 194
rect 152 185 157 194
rect 143 179 157 185
rect 143 170 148 179
rect 152 170 157 179
rect 143 164 157 170
rect 143 155 148 164
rect 152 155 157 164
rect 143 144 157 155
rect 143 140 148 144
rect 152 140 157 144
rect 143 134 157 140
rect 143 125 148 134
rect 152 125 157 134
rect 143 119 157 125
rect 143 110 148 119
rect 152 110 157 119
rect 143 104 157 110
rect 143 95 148 104
rect 152 95 157 104
rect 143 89 157 95
rect 143 85 148 89
rect 152 85 157 89
rect 143 74 157 85
rect 143 65 148 74
rect 152 65 157 74
rect 143 59 157 65
rect 143 55 148 59
rect 152 55 157 59
rect 14 31 30 33
rect 14 29 39 31
rect 14 25 17 29
rect 21 25 23 29
rect 37 27 39 29
rect 43 27 53 32
rect 37 25 53 27
rect 14 19 53 25
rect 14 15 23 19
rect 37 18 53 19
rect 57 31 138 32
rect 57 18 64 31
rect 37 17 64 18
rect 68 17 74 31
rect 78 17 84 31
rect 88 17 94 31
rect 98 17 104 31
rect 108 17 114 31
rect 118 30 138 31
rect 143 30 157 55
rect 162 31 262 32
rect 162 30 182 31
rect 118 17 182 30
rect 186 17 192 31
rect 196 17 202 31
rect 206 17 212 31
rect 216 17 222 31
rect 226 17 232 31
rect 236 17 242 31
rect 246 30 262 31
rect 270 30 276 229
rect 246 17 263 30
rect 37 16 263 17
rect 267 16 276 30
rect 37 15 276 16
rect 14 14 276 15
rect 280 14 281 243
<< nsubstratendiff >>
rect 19 647 281 648
rect 19 645 148 647
rect 19 640 45 645
rect 19 626 20 640
rect 29 636 45 640
rect 54 636 56 645
rect 60 636 66 645
rect 75 636 81 645
rect 90 636 96 645
rect 105 636 111 645
rect 115 643 148 645
rect 152 645 281 647
rect 152 643 183 645
rect 115 637 183 643
rect 115 636 148 637
rect 29 630 36 636
rect 140 630 148 636
rect 29 626 30 630
rect 141 629 148 630
rect 19 620 30 626
rect 19 606 20 620
rect 29 606 30 620
rect 19 600 30 606
rect 19 586 20 600
rect 29 586 30 600
rect 19 580 30 586
rect 19 566 20 580
rect 29 566 30 580
rect 19 560 30 566
rect 19 546 20 560
rect 29 546 30 560
rect 19 540 30 546
rect 19 526 20 540
rect 29 526 30 540
rect 19 520 30 526
rect 19 506 20 520
rect 29 506 30 520
rect 19 500 30 506
rect 19 486 20 500
rect 29 486 30 500
rect 19 480 30 486
rect 19 466 20 480
rect 29 466 30 480
rect 19 460 30 466
rect 19 446 20 460
rect 29 446 30 460
rect 142 623 148 629
rect 152 636 183 637
rect 187 636 193 645
rect 202 636 208 645
rect 217 636 223 645
rect 232 636 238 645
rect 242 636 244 645
rect 253 640 281 645
rect 253 636 271 640
rect 152 630 160 636
rect 264 630 271 636
rect 152 629 159 630
rect 152 623 158 629
rect 142 617 158 623
rect 142 603 148 617
rect 152 603 158 617
rect 142 597 158 603
rect 142 583 148 597
rect 152 583 158 597
rect 142 577 158 583
rect 142 563 148 577
rect 152 563 158 577
rect 142 557 158 563
rect 142 543 148 557
rect 152 543 158 557
rect 142 537 158 543
rect 142 523 148 537
rect 152 523 158 537
rect 142 517 158 523
rect 142 503 148 517
rect 152 503 158 517
rect 142 497 158 503
rect 142 483 148 497
rect 152 483 158 497
rect 142 477 158 483
rect 142 463 148 477
rect 152 463 158 477
rect 142 457 158 463
rect 19 440 30 446
rect 38 441 138 442
rect 38 440 51 441
rect 19 431 20 440
rect 29 437 51 440
rect 55 437 61 441
rect 70 437 76 441
rect 85 437 91 441
rect 100 437 106 441
rect 115 440 138 441
rect 142 443 148 457
rect 152 443 158 457
rect 270 626 271 630
rect 280 626 281 640
rect 270 620 281 626
rect 270 606 271 620
rect 280 606 281 620
rect 270 600 281 606
rect 270 586 271 600
rect 280 586 281 600
rect 270 580 281 586
rect 270 566 271 580
rect 280 566 281 580
rect 270 560 281 566
rect 270 546 271 560
rect 280 546 281 560
rect 270 540 281 546
rect 270 526 271 540
rect 280 526 281 540
rect 270 520 281 526
rect 270 506 271 520
rect 280 506 281 520
rect 270 500 281 506
rect 270 486 271 500
rect 280 486 281 500
rect 270 480 281 486
rect 270 466 271 480
rect 280 466 281 480
rect 270 460 281 466
rect 142 440 158 443
rect 162 441 262 442
rect 162 440 184 441
rect 115 437 184 440
rect 193 437 199 441
rect 208 437 214 441
rect 223 437 229 441
rect 238 437 244 441
rect 248 440 262 441
rect 270 446 271 460
rect 280 446 281 460
rect 270 440 281 446
rect 248 437 271 440
rect 29 435 148 437
rect 29 431 46 435
rect 115 433 148 435
rect 152 435 271 437
rect 152 433 184 435
rect 115 431 184 433
rect 253 431 271 435
rect 280 431 281 440
rect 19 430 281 431
rect 0 331 295 332
rect 0 2 2 331
rect 6 329 17 331
rect 6 326 7 329
rect 15 327 17 329
rect 21 329 38 331
rect 21 327 23 329
rect 15 326 23 327
rect 31 327 38 329
rect 42 327 45 331
rect 49 329 64 331
rect 49 327 50 329
rect 31 326 50 327
rect 63 327 64 329
rect 68 327 74 331
rect 83 329 98 331
rect 83 327 84 329
rect 63 326 84 327
rect 63 324 67 326
rect 79 324 83 326
rect 97 327 98 329
rect 102 327 109 331
rect 113 329 137 331
rect 113 327 122 329
rect 97 326 122 327
rect 111 324 115 326
rect 135 327 137 329
rect 141 327 194 331
rect 203 327 209 331
rect 213 327 223 331
rect 227 329 242 331
rect 227 327 228 329
rect 135 326 228 327
rect 192 324 197 326
rect 209 324 213 326
rect 225 324 228 326
rect 241 327 242 329
rect 251 327 257 331
rect 261 327 271 331
rect 275 329 295 331
rect 275 327 276 329
rect 241 326 276 327
rect 241 324 245 326
rect 257 324 261 326
rect 273 324 276 326
rect 289 324 295 329
rect 293 323 295 324
rect 299 323 300 332
rect 36 261 43 265
rect 79 265 83 266
rect 192 265 197 266
rect 241 265 245 266
rect 56 264 241 265
rect 56 263 193 264
rect 56 261 59 263
rect 6 259 59 261
rect 113 260 193 263
rect 197 261 241 264
rect 245 261 289 265
rect 197 260 289 261
rect 113 259 263 260
rect 6 258 240 259
rect 6 254 17 258
rect 36 257 194 258
rect 36 254 54 257
rect 6 253 54 254
rect 108 254 194 257
rect 228 255 240 258
rect 254 256 263 259
rect 287 257 289 260
rect 293 257 300 323
rect 287 256 300 257
rect 254 255 300 256
rect 228 254 300 255
rect 108 253 300 254
rect 6 252 300 253
rect 6 8 8 252
rect 289 251 300 252
rect 289 8 290 251
rect 6 6 290 8
rect 6 2 8 6
rect 287 2 290 6
rect 299 2 300 251
rect 0 0 300 2
<< psubstratepcontact >>
rect 1 658 115 667
rect 184 658 298 667
rect 1 415 10 654
rect 15 410 29 419
rect 39 410 113 419
rect 148 410 152 419
rect 184 410 288 419
rect 290 412 299 656
rect 1 343 5 407
rect 295 402 299 406
rect 295 392 299 396
rect 295 382 299 386
rect 295 372 299 376
rect 295 362 299 366
rect 17 343 21 347
rect 38 342 42 346
rect 45 342 49 346
rect 64 342 83 346
rect 99 343 103 347
rect 108 343 112 347
rect 124 343 128 347
rect 194 342 213 346
rect 223 343 227 347
rect 295 352 299 356
rect 242 342 251 346
rect 257 342 261 346
rect 271 342 275 346
rect 290 342 299 346
rect 17 236 36 240
rect 53 237 117 241
rect 17 228 26 232
rect 17 208 26 222
rect 54 229 63 233
rect 69 229 78 233
rect 84 229 93 233
rect 99 229 108 233
rect 114 229 118 233
rect 148 230 152 239
rect 182 237 246 241
rect 17 188 26 202
rect 17 168 26 182
rect 17 148 26 162
rect 17 128 26 142
rect 17 108 26 122
rect 17 88 26 102
rect 17 68 26 82
rect 17 48 26 62
rect 17 33 26 42
rect 148 215 152 224
rect 182 229 191 233
rect 197 229 206 233
rect 212 229 221 233
rect 227 229 236 233
rect 242 229 246 233
rect 270 229 274 243
rect 148 200 152 209
rect 148 185 152 194
rect 148 170 152 179
rect 148 155 152 164
rect 148 140 152 144
rect 148 125 152 134
rect 148 110 152 119
rect 148 95 152 104
rect 148 85 152 89
rect 148 65 152 74
rect 148 55 152 59
rect 17 25 21 29
rect 23 25 37 29
rect 39 27 43 31
rect 23 15 37 19
rect 53 18 57 32
rect 64 17 68 31
rect 74 17 78 31
rect 84 17 88 31
rect 94 17 98 31
rect 104 17 108 31
rect 114 17 118 31
rect 182 17 186 31
rect 192 17 196 31
rect 202 17 206 31
rect 212 17 216 31
rect 222 17 226 31
rect 232 17 236 31
rect 242 17 246 31
rect 263 16 267 30
rect 276 14 280 243
<< nsubstratencontact >>
rect 20 626 29 640
rect 45 636 54 645
rect 56 636 60 645
rect 66 636 75 645
rect 81 636 90 645
rect 96 636 105 645
rect 111 636 115 645
rect 148 643 152 647
rect 20 606 29 620
rect 20 586 29 600
rect 20 566 29 580
rect 20 546 29 560
rect 20 526 29 540
rect 20 506 29 520
rect 20 486 29 500
rect 20 466 29 480
rect 20 446 29 460
rect 148 623 152 637
rect 183 636 187 645
rect 193 636 202 645
rect 208 636 217 645
rect 223 636 232 645
rect 238 636 242 645
rect 244 636 253 645
rect 148 603 152 617
rect 148 583 152 597
rect 148 563 152 577
rect 148 543 152 557
rect 148 523 152 537
rect 148 503 152 517
rect 148 483 152 497
rect 148 463 152 477
rect 20 431 29 440
rect 51 437 55 441
rect 61 437 70 441
rect 76 437 85 441
rect 91 437 100 441
rect 106 437 115 441
rect 148 443 152 457
rect 271 626 280 640
rect 271 606 280 620
rect 271 586 280 600
rect 271 566 280 580
rect 271 546 280 560
rect 271 526 280 540
rect 271 506 280 520
rect 271 486 280 500
rect 271 466 280 480
rect 184 437 193 441
rect 199 437 208 441
rect 214 437 223 441
rect 229 437 238 441
rect 244 437 248 441
rect 271 446 280 460
rect 46 431 115 435
rect 148 433 152 437
rect 184 431 253 435
rect 271 431 280 440
rect 2 2 6 331
rect 17 327 21 331
rect 38 327 42 331
rect 45 327 49 331
rect 64 327 68 331
rect 74 327 83 331
rect 98 327 102 331
rect 109 327 113 331
rect 137 327 141 331
rect 194 327 203 331
rect 209 327 213 331
rect 223 327 227 331
rect 242 327 251 331
rect 257 327 261 331
rect 271 327 275 331
rect 295 323 299 332
rect 59 259 113 263
rect 193 260 197 264
rect 241 261 245 265
rect 17 254 36 258
rect 54 253 108 257
rect 194 254 228 258
rect 240 255 254 259
rect 263 256 287 260
rect 8 2 287 6
rect 290 2 299 251
<< polysilicon >>
rect 31 624 38 627
rect 138 624 141 627
rect 31 614 37 624
rect 31 595 32 614
rect 36 595 37 614
rect 31 583 37 595
rect 139 583 141 624
rect 31 580 38 583
rect 138 580 141 583
rect 31 562 37 580
rect 139 562 141 580
rect 31 559 38 562
rect 138 559 141 562
rect 31 549 37 559
rect 31 530 32 549
rect 36 530 37 549
rect 31 519 37 530
rect 139 519 141 559
rect 31 516 38 519
rect 138 516 141 519
rect 31 498 37 516
rect 139 498 141 516
rect 31 495 38 498
rect 138 495 141 498
rect 31 481 37 495
rect 31 452 32 481
rect 36 454 37 481
rect 139 454 141 495
rect 36 452 38 454
rect 31 451 38 452
rect 138 451 141 454
rect 159 624 162 627
rect 262 624 269 627
rect 159 583 161 624
rect 263 612 269 624
rect 263 593 264 612
rect 268 593 269 612
rect 263 583 269 593
rect 159 580 162 583
rect 262 580 269 583
rect 159 562 161 580
rect 263 562 269 580
rect 159 559 162 562
rect 262 559 269 562
rect 159 519 161 559
rect 263 549 269 559
rect 263 530 264 549
rect 268 530 269 549
rect 263 519 269 530
rect 159 516 162 519
rect 262 516 269 519
rect 159 498 161 516
rect 263 498 269 516
rect 159 495 162 498
rect 262 495 269 498
rect 159 454 161 495
rect 263 484 269 495
rect 263 455 264 484
rect 268 455 269 484
rect 263 454 269 455
rect 159 451 162 454
rect 262 451 269 454
rect 111 404 126 405
rect 125 395 126 404
rect 191 399 210 405
rect 191 395 193 399
rect 207 395 210 399
rect 274 404 290 405
rect 274 395 275 404
rect 289 395 290 404
rect 207 390 208 395
rect 24 389 35 390
rect 24 385 25 389
rect 34 385 35 389
rect 19 383 21 385
rect 24 384 35 385
rect 44 384 78 386
rect 27 383 29 384
rect 44 383 46 384
rect 52 383 54 384
rect 60 383 62 384
rect 68 383 70 384
rect 76 383 78 384
rect 84 384 118 386
rect 84 383 86 384
rect 92 383 94 384
rect 100 383 102 384
rect 108 383 110 384
rect 116 383 118 384
rect 124 383 126 385
rect 132 383 134 385
rect 140 383 142 385
rect 148 383 150 385
rect 198 383 200 390
rect 206 384 216 386
rect 206 383 208 384
rect 214 383 216 384
rect 222 384 232 386
rect 222 383 224 384
rect 230 383 232 384
rect 238 383 240 385
rect 246 383 248 385
rect 254 384 264 386
rect 254 383 256 384
rect 262 383 264 384
rect 270 384 280 386
rect 270 383 272 384
rect 278 383 280 384
rect 286 383 288 386
rect 19 352 21 353
rect 27 352 29 353
rect 8 351 21 352
rect 8 347 9 351
rect 13 350 21 351
rect 24 351 30 352
rect 13 347 14 350
rect 8 346 14 347
rect 24 347 25 351
rect 29 347 30 351
rect 44 350 46 353
rect 52 351 54 353
rect 60 351 62 353
rect 24 346 30 347
rect 51 350 62 351
rect 51 346 52 350
rect 61 346 62 350
rect 51 345 62 346
rect 68 350 70 353
rect 76 350 78 353
rect 84 352 86 353
rect 92 352 94 353
rect 84 351 96 352
rect 84 349 86 351
rect 85 347 86 349
rect 95 347 96 351
rect 100 350 102 353
rect 108 350 110 353
rect 116 350 118 353
rect 124 352 126 353
rect 132 352 134 353
rect 140 352 142 353
rect 148 352 150 353
rect 124 351 150 352
rect 124 350 137 351
rect 85 346 96 347
rect 136 347 137 350
rect 146 350 150 351
rect 198 352 200 353
rect 206 352 208 353
rect 198 350 208 352
rect 214 352 216 353
rect 222 352 224 353
rect 214 350 224 352
rect 230 352 232 353
rect 238 352 240 353
rect 146 347 147 350
rect 136 346 147 347
rect 229 351 240 352
rect 229 347 230 351
rect 239 347 240 351
rect 229 346 240 347
rect 246 352 248 353
rect 254 352 256 353
rect 246 350 256 352
rect 262 352 264 353
rect 270 352 272 353
rect 262 350 272 352
rect 278 352 280 353
rect 286 352 288 353
rect 277 351 288 352
rect 277 347 278 351
rect 287 347 288 351
rect 277 346 288 347
rect 31 339 147 340
rect 31 335 32 339
rect 41 335 80 339
rect 89 335 137 339
rect 146 335 147 339
rect 31 334 147 335
rect 8 327 14 328
rect 8 323 9 327
rect 13 324 14 327
rect 24 327 30 328
rect 13 323 21 324
rect 8 322 21 323
rect 24 323 25 327
rect 29 323 30 327
rect 51 327 62 328
rect 51 323 52 327
rect 61 323 62 327
rect 24 322 30 323
rect 19 321 21 322
rect 27 321 29 322
rect 44 321 46 323
rect 51 322 62 323
rect 52 321 54 322
rect 60 321 62 322
rect 85 327 96 328
rect 85 324 86 327
rect 68 321 70 323
rect 76 321 78 323
rect 84 323 86 324
rect 95 323 96 327
rect 123 327 134 328
rect 84 322 96 323
rect 84 321 86 322
rect 92 321 94 322
rect 100 321 102 323
rect 108 321 110 323
rect 123 323 124 327
rect 133 324 134 327
rect 133 323 150 324
rect 116 321 118 323
rect 123 322 150 323
rect 124 321 126 322
rect 132 321 134 322
rect 140 321 142 322
rect 148 321 150 322
rect 198 323 208 325
rect 198 321 200 323
rect 206 321 208 323
rect 214 323 224 325
rect 214 321 216 323
rect 222 321 224 323
rect 229 327 240 328
rect 229 323 230 327
rect 239 323 240 327
rect 229 322 240 323
rect 230 321 232 322
rect 238 321 240 322
rect 246 322 256 324
rect 246 321 248 322
rect 254 321 256 322
rect 262 322 272 324
rect 262 321 264 322
rect 270 321 272 322
rect 277 327 288 328
rect 277 323 278 327
rect 287 323 288 327
rect 277 322 288 323
rect 278 321 280 322
rect 286 321 288 322
rect 19 268 21 269
rect 27 268 29 269
rect 44 268 46 269
rect 52 268 54 269
rect 60 268 62 269
rect 68 268 70 269
rect 76 268 78 269
rect 10 267 21 268
rect 10 263 11 267
rect 20 263 21 267
rect 10 262 21 263
rect 24 267 35 268
rect 24 263 25 267
rect 34 263 35 267
rect 44 267 78 268
rect 24 262 35 263
rect 44 263 45 267
rect 54 266 78 267
rect 84 268 86 269
rect 92 268 94 269
rect 100 268 102 269
rect 108 268 110 269
rect 116 268 118 269
rect 84 266 118 268
rect 124 267 126 269
rect 132 267 134 269
rect 140 267 142 269
rect 148 267 150 269
rect 198 267 200 269
rect 206 268 208 269
rect 214 268 216 269
rect 206 266 216 268
rect 222 268 224 269
rect 230 268 232 269
rect 222 266 232 268
rect 238 267 240 269
rect 246 267 248 269
rect 254 268 256 269
rect 262 268 264 269
rect 254 266 264 268
rect 270 268 272 269
rect 278 268 280 269
rect 270 266 280 268
rect 286 267 288 269
rect 54 263 55 266
rect 44 262 55 263
rect 31 217 38 219
rect 31 43 32 217
rect 36 216 38 217
rect 138 216 142 219
rect 36 174 37 216
rect 139 174 142 216
rect 36 171 38 174
rect 138 171 142 174
rect 36 153 37 171
rect 139 153 142 171
rect 36 150 38 153
rect 138 150 142 153
rect 36 109 37 150
rect 139 109 142 150
rect 36 106 38 109
rect 138 106 142 109
rect 36 88 37 106
rect 139 88 142 106
rect 36 85 38 88
rect 138 85 142 88
rect 36 44 37 85
rect 139 44 142 85
rect 36 43 38 44
rect 31 41 38 43
rect 138 41 142 44
rect 158 216 162 219
rect 262 217 269 219
rect 262 216 264 217
rect 158 174 161 216
rect 263 174 264 216
rect 158 171 162 174
rect 262 171 264 174
rect 158 153 161 171
rect 263 153 264 171
rect 158 150 162 153
rect 262 150 264 153
rect 158 109 161 150
rect 263 109 264 150
rect 158 106 162 109
rect 262 106 264 109
rect 158 88 161 106
rect 263 88 264 106
rect 158 85 162 88
rect 262 85 264 88
rect 158 44 161 85
rect 263 44 264 85
rect 158 41 162 44
rect 262 43 264 44
rect 268 43 269 217
rect 262 41 269 43
<< polycontact >>
rect 32 595 36 614
rect 32 530 36 549
rect 32 452 36 481
rect 264 593 268 612
rect 264 530 268 549
rect 264 455 268 484
rect 111 395 125 404
rect 193 390 207 399
rect 275 395 289 404
rect 25 385 34 389
rect 9 347 13 351
rect 25 347 29 351
rect 52 346 61 350
rect 86 347 95 351
rect 137 347 146 351
rect 230 347 239 351
rect 278 347 287 351
rect 32 335 41 339
rect 80 335 89 339
rect 137 335 146 339
rect 9 323 13 327
rect 25 323 29 327
rect 52 323 61 327
rect 86 323 95 327
rect 124 323 133 327
rect 230 323 239 327
rect 278 323 287 327
rect 11 263 20 267
rect 25 263 34 267
rect 45 263 54 267
rect 32 43 36 217
rect 264 43 268 217
<< metal1 >>
rect 20 997 280 1000
rect 20 743 23 997
rect 277 743 280 997
rect 20 740 280 743
rect 62 700 238 740
rect 102 690 198 700
rect 112 680 188 690
rect 0 667 116 669
rect 0 658 1 667
rect 115 658 116 667
rect 0 654 10 658
rect 0 415 1 654
rect 14 654 117 655
rect 18 650 22 654
rect 111 650 117 654
rect 18 645 117 650
rect 18 641 22 645
rect 26 641 30 645
rect 18 640 30 641
rect 18 626 20 640
rect 29 631 30 640
rect 44 636 45 645
rect 54 636 56 645
rect 60 636 61 645
rect 44 634 61 636
rect 44 631 45 634
rect 29 630 45 631
rect 54 630 56 634
rect 60 631 61 634
rect 65 636 66 645
rect 75 636 76 645
rect 65 634 76 636
rect 65 631 66 634
rect 60 630 66 631
rect 75 631 76 634
rect 80 636 81 645
rect 90 636 91 645
rect 80 634 91 636
rect 80 631 81 634
rect 75 630 81 631
rect 90 631 91 634
rect 95 636 96 645
rect 105 636 106 645
rect 95 634 106 636
rect 95 631 96 634
rect 90 630 96 631
rect 105 631 106 634
rect 110 636 111 645
rect 115 636 117 645
rect 110 634 117 636
rect 110 631 111 634
rect 105 630 111 631
rect 115 630 117 634
rect 29 626 117 630
rect 18 625 117 626
rect 18 621 20 625
rect 29 621 32 625
rect 36 622 117 625
rect 36 621 52 622
rect 18 620 41 621
rect 18 606 20 620
rect 29 617 41 620
rect 18 605 29 606
rect 18 601 20 605
rect 18 600 29 601
rect 18 586 20 600
rect 39 592 41 617
rect 29 589 41 592
rect 29 586 32 589
rect 18 585 32 586
rect 18 581 20 585
rect 29 581 32 585
rect 18 580 32 581
rect 18 566 20 580
rect 29 566 32 580
rect 18 565 32 566
rect 18 561 20 565
rect 29 561 32 565
rect 18 560 32 561
rect 18 546 20 560
rect 29 555 32 560
rect 36 587 41 589
rect 50 618 52 621
rect 116 618 117 622
rect 50 617 117 618
rect 120 654 180 680
rect 184 667 300 669
rect 298 658 300 667
rect 290 656 300 658
rect 50 592 52 617
rect 120 612 143 654
rect 56 608 143 612
rect 120 599 143 608
rect 56 595 143 599
rect 50 590 117 592
rect 50 587 52 590
rect 36 586 52 587
rect 116 586 117 590
rect 36 576 117 586
rect 36 572 41 576
rect 60 572 61 576
rect 70 572 71 576
rect 75 572 76 576
rect 85 572 86 576
rect 90 572 91 576
rect 100 572 101 576
rect 105 572 106 576
rect 115 572 117 576
rect 36 570 117 572
rect 36 566 41 570
rect 60 566 61 570
rect 70 566 71 570
rect 75 566 76 570
rect 85 566 86 570
rect 90 566 91 570
rect 100 566 101 570
rect 105 566 106 570
rect 115 566 117 570
rect 36 556 117 566
rect 36 555 42 556
rect 29 552 42 555
rect 18 545 29 546
rect 18 541 20 545
rect 18 540 29 541
rect 18 526 20 540
rect 39 527 42 552
rect 29 526 42 527
rect 18 525 42 526
rect 18 521 20 525
rect 29 524 42 525
rect 29 521 32 524
rect 18 520 32 521
rect 18 506 20 520
rect 29 506 32 520
rect 18 505 32 506
rect 18 501 20 505
rect 29 501 32 505
rect 18 500 32 501
rect 18 486 20 500
rect 29 490 32 500
rect 36 522 42 524
rect 51 552 55 556
rect 114 552 117 556
rect 51 527 52 552
rect 120 548 143 595
rect 55 543 143 548
rect 55 534 56 543
rect 120 534 143 543
rect 55 530 143 534
rect 51 526 117 527
rect 51 522 55 526
rect 114 522 117 526
rect 36 512 117 522
rect 36 508 41 512
rect 60 508 61 512
rect 70 508 71 512
rect 75 508 76 512
rect 85 508 86 512
rect 90 508 91 512
rect 100 508 101 512
rect 105 508 106 512
rect 115 508 117 512
rect 36 506 117 508
rect 36 502 41 506
rect 60 502 61 506
rect 70 502 71 506
rect 75 502 76 506
rect 85 502 86 506
rect 90 502 91 506
rect 100 502 101 506
rect 105 502 106 506
rect 115 502 117 506
rect 36 493 117 502
rect 36 492 55 493
rect 36 490 42 492
rect 29 488 42 490
rect 18 485 29 486
rect 18 481 20 485
rect 18 480 29 481
rect 18 466 20 480
rect 18 465 29 466
rect 18 461 20 465
rect 18 460 29 461
rect 18 446 20 460
rect 18 445 29 446
rect 18 441 20 445
rect 18 440 29 441
rect 14 431 20 440
rect 14 430 29 431
rect 32 436 36 452
rect 39 458 42 488
rect 51 489 55 492
rect 114 489 117 493
rect 51 488 117 489
rect 51 462 52 488
rect 120 483 143 530
rect 55 479 143 483
rect 55 470 56 479
rect 120 470 143 479
rect 55 466 143 470
rect 51 461 116 462
rect 51 458 54 461
rect 39 457 54 458
rect 113 457 116 461
rect 39 447 116 457
rect 39 443 40 447
rect 49 443 51 447
rect 60 443 61 447
rect 70 443 71 447
rect 75 443 76 447
rect 85 443 86 447
rect 90 443 91 447
rect 100 443 101 447
rect 105 443 106 447
rect 115 443 116 447
rect 39 441 116 443
rect 39 439 46 441
rect 44 437 46 439
rect 50 437 51 441
rect 55 437 56 441
rect 60 437 61 441
rect 70 437 71 441
rect 75 437 76 441
rect 85 437 86 441
rect 90 437 91 441
rect 100 437 101 441
rect 105 437 106 441
rect 115 437 116 441
rect 32 435 41 436
rect 32 430 41 431
rect 44 435 116 437
rect 44 431 46 435
rect 115 431 116 435
rect 44 430 116 431
rect 10 421 15 425
rect 10 419 29 421
rect 10 415 15 419
rect 0 410 15 415
rect 0 409 29 410
rect 0 407 7 409
rect 0 343 1 407
rect 5 395 7 407
rect 11 405 13 409
rect 27 405 29 409
rect 11 404 29 405
rect 5 393 11 395
rect 32 398 36 430
rect 113 421 115 425
rect 39 419 115 421
rect 113 410 115 419
rect 39 409 108 410
rect 120 407 143 466
rect 147 647 153 648
rect 147 643 148 647
rect 152 643 153 647
rect 147 642 153 643
rect 147 638 148 642
rect 152 638 153 642
rect 147 637 153 638
rect 147 623 148 637
rect 152 623 153 637
rect 147 622 153 623
rect 147 618 148 622
rect 152 618 153 622
rect 147 617 153 618
rect 147 603 148 617
rect 152 603 153 617
rect 147 602 153 603
rect 147 598 148 602
rect 152 598 153 602
rect 147 597 153 598
rect 147 583 148 597
rect 152 583 153 597
rect 147 582 153 583
rect 147 578 148 582
rect 152 578 153 582
rect 147 577 153 578
rect 147 563 148 577
rect 152 563 153 577
rect 147 562 153 563
rect 147 558 148 562
rect 152 558 153 562
rect 147 557 153 558
rect 147 543 148 557
rect 152 543 153 557
rect 147 542 153 543
rect 147 538 148 542
rect 152 538 153 542
rect 147 537 153 538
rect 147 523 148 537
rect 152 523 153 537
rect 147 522 153 523
rect 147 518 148 522
rect 152 518 153 522
rect 147 517 153 518
rect 147 503 148 517
rect 152 503 153 517
rect 147 502 153 503
rect 147 498 148 502
rect 152 498 153 502
rect 147 497 153 498
rect 147 483 148 497
rect 152 483 153 497
rect 147 482 153 483
rect 147 478 148 482
rect 152 478 153 482
rect 147 477 153 478
rect 147 463 148 477
rect 152 463 153 477
rect 147 462 153 463
rect 147 458 148 462
rect 152 458 153 462
rect 147 457 153 458
rect 147 443 148 457
rect 152 443 153 457
rect 147 442 153 443
rect 147 438 148 442
rect 152 438 153 442
rect 147 437 153 438
rect 147 433 148 437
rect 152 433 153 437
rect 147 430 153 433
rect 157 612 180 654
rect 183 651 189 655
rect 278 651 282 655
rect 183 645 282 651
rect 187 636 188 645
rect 183 634 188 636
rect 187 631 188 634
rect 192 636 193 645
rect 202 636 203 645
rect 192 634 203 636
rect 192 631 193 634
rect 187 630 193 631
rect 202 631 203 634
rect 207 636 208 645
rect 217 636 218 645
rect 207 634 218 636
rect 207 631 208 634
rect 202 630 208 631
rect 217 631 218 634
rect 222 636 223 645
rect 232 636 233 645
rect 222 634 233 636
rect 222 631 223 634
rect 217 630 223 631
rect 232 631 233 634
rect 237 636 238 645
rect 242 636 244 645
rect 253 636 254 645
rect 237 634 254 636
rect 237 631 238 634
rect 232 630 238 631
rect 242 630 244 634
rect 253 631 254 634
rect 268 641 271 645
rect 280 641 282 645
rect 268 640 282 641
rect 268 631 271 640
rect 253 630 271 631
rect 183 626 271 630
rect 280 626 282 640
rect 183 625 282 626
rect 183 622 264 625
rect 183 618 186 622
rect 245 621 264 622
rect 268 621 271 625
rect 280 621 282 625
rect 245 620 282 621
rect 245 618 249 620
rect 183 616 249 618
rect 157 608 244 612
rect 157 599 180 608
rect 157 595 244 599
rect 157 548 180 595
rect 248 590 249 616
rect 183 589 249 590
rect 183 585 186 589
rect 245 586 249 589
rect 258 616 271 620
rect 258 590 261 616
rect 280 606 282 620
rect 271 605 282 606
rect 280 601 282 605
rect 271 600 282 601
rect 258 588 271 590
rect 258 586 264 588
rect 245 585 264 586
rect 183 576 264 585
rect 183 572 184 576
rect 193 572 194 576
rect 198 572 199 576
rect 208 572 209 576
rect 213 572 214 576
rect 223 572 224 576
rect 228 572 229 576
rect 238 572 239 576
rect 258 572 264 576
rect 183 570 264 572
rect 183 566 184 570
rect 193 566 194 570
rect 198 566 199 570
rect 208 566 209 570
rect 213 566 214 570
rect 223 566 224 570
rect 228 566 229 570
rect 238 566 239 570
rect 258 566 264 570
rect 183 557 264 566
rect 183 553 186 557
rect 245 556 264 557
rect 245 553 249 556
rect 183 552 249 553
rect 157 543 244 548
rect 157 534 180 543
rect 157 530 244 534
rect 157 483 180 530
rect 248 527 249 552
rect 183 526 249 527
rect 183 522 186 526
rect 245 522 249 526
rect 258 554 264 556
rect 268 586 271 588
rect 280 586 282 600
rect 268 585 282 586
rect 268 581 271 585
rect 280 581 282 585
rect 268 580 282 581
rect 268 566 271 580
rect 280 566 282 580
rect 268 565 282 566
rect 268 561 271 565
rect 280 561 282 565
rect 268 560 282 561
rect 268 554 271 560
rect 258 552 271 554
rect 258 527 261 552
rect 280 546 282 560
rect 271 545 282 546
rect 280 541 282 545
rect 271 540 282 541
rect 258 526 271 527
rect 280 526 282 540
rect 258 525 282 526
rect 258 524 271 525
rect 258 522 264 524
rect 183 512 264 522
rect 192 508 193 512
rect 197 508 198 512
rect 207 508 208 512
rect 212 508 213 512
rect 222 508 223 512
rect 227 508 228 512
rect 237 508 238 512
rect 257 508 264 512
rect 183 506 264 508
rect 192 502 193 506
rect 197 502 198 506
rect 207 502 208 506
rect 212 502 213 506
rect 222 502 223 506
rect 227 502 228 506
rect 237 502 238 506
rect 257 502 264 506
rect 183 493 264 502
rect 183 489 184 493
rect 248 492 264 493
rect 248 489 250 492
rect 183 488 250 489
rect 157 479 244 483
rect 157 470 180 479
rect 157 466 244 470
rect 148 419 152 421
rect 157 407 180 466
rect 248 462 250 488
rect 184 461 250 462
rect 184 457 187 461
rect 246 458 250 461
rect 259 490 264 492
rect 268 521 271 524
rect 280 521 282 525
rect 268 520 282 521
rect 268 506 271 520
rect 280 506 282 520
rect 268 505 282 506
rect 268 501 271 505
rect 280 501 282 505
rect 268 500 282 501
rect 268 490 271 500
rect 259 488 271 490
rect 259 458 261 488
rect 280 486 282 500
rect 271 485 282 486
rect 246 457 261 458
rect 184 447 261 457
rect 193 443 194 447
rect 198 443 199 447
rect 208 443 209 447
rect 213 443 214 447
rect 223 443 224 447
rect 228 443 229 447
rect 238 443 239 447
rect 243 443 245 447
rect 254 443 256 447
rect 260 443 261 447
rect 184 441 261 443
rect 193 437 194 441
rect 198 437 199 441
rect 208 437 209 441
rect 213 437 214 441
rect 223 437 224 441
rect 228 437 229 441
rect 238 437 239 441
rect 243 437 244 441
rect 248 437 249 441
rect 253 439 261 441
rect 253 437 256 439
rect 184 435 256 437
rect 264 436 268 455
rect 253 431 256 435
rect 184 430 256 431
rect 259 435 268 436
rect 259 430 268 431
rect 280 481 282 485
rect 271 480 282 481
rect 280 466 282 480
rect 271 465 282 466
rect 280 461 282 465
rect 271 460 282 461
rect 280 446 282 460
rect 271 445 282 446
rect 280 441 282 445
rect 271 440 286 441
rect 280 431 286 440
rect 271 430 286 431
rect 288 421 290 425
rect 184 419 290 421
rect 288 412 290 419
rect 299 412 300 656
rect 288 411 300 412
rect 288 410 295 411
rect 293 407 295 410
rect 299 407 300 411
rect 39 404 108 405
rect 111 404 290 407
rect 32 393 41 398
rect 125 403 275 404
rect 125 395 190 403
rect 111 393 190 395
rect 5 354 7 393
rect 37 390 41 393
rect 14 385 25 389
rect 37 387 131 390
rect 134 388 190 393
rect 193 399 208 400
rect 207 390 208 399
rect 211 395 275 403
rect 289 395 290 404
rect 293 406 300 407
rect 293 402 295 406
rect 299 402 300 406
rect 293 401 300 402
rect 293 397 295 401
rect 299 397 300 401
rect 293 396 300 397
rect 211 390 228 395
rect 293 392 295 396
rect 299 392 300 396
rect 127 385 131 387
rect 150 387 190 388
rect 211 387 215 390
rect 150 385 215 387
rect 293 391 300 392
rect 293 388 295 391
rect 289 387 295 388
rect 299 387 300 391
rect 289 386 300 387
rect 14 380 18 385
rect 14 360 18 361
rect 22 380 26 382
rect 22 375 26 376
rect 22 370 26 371
rect 22 365 26 366
rect 22 360 26 361
rect 19 356 22 357
rect 19 354 26 356
rect 30 379 34 382
rect 39 381 123 384
rect 39 379 43 381
rect 55 379 59 381
rect 47 373 51 374
rect 47 368 51 369
rect 47 363 51 364
rect 47 358 51 359
rect 34 355 35 358
rect 30 354 35 355
rect 5 343 6 354
rect 0 341 6 343
rect 19 348 22 354
rect 16 347 22 348
rect 0 331 6 332
rect 0 2 2 331
rect 9 327 12 347
rect 16 343 17 347
rect 21 343 22 347
rect 16 342 22 343
rect 25 339 28 347
rect 32 339 35 354
rect 38 354 47 357
rect 71 379 75 381
rect 63 373 67 374
rect 63 368 67 369
rect 63 363 67 364
rect 63 358 67 359
rect 87 379 91 381
rect 79 373 83 374
rect 79 368 83 369
rect 79 363 83 364
rect 79 358 83 359
rect 38 346 49 354
rect 64 352 67 354
rect 103 380 107 381
rect 95 373 99 374
rect 95 368 99 369
rect 95 363 99 364
rect 95 358 99 359
rect 119 379 123 381
rect 111 373 115 374
rect 111 368 115 369
rect 111 363 115 364
rect 119 364 123 365
rect 127 382 147 385
rect 158 383 215 385
rect 218 383 237 386
rect 127 378 131 382
rect 143 379 147 382
rect 111 358 115 359
rect 79 352 83 354
rect 64 346 83 352
rect 111 348 115 354
rect 42 342 45 346
rect 16 331 22 332
rect 16 327 17 331
rect 21 327 22 331
rect 16 326 22 327
rect 6 318 11 320
rect 6 274 7 318
rect 19 317 22 326
rect 25 327 28 335
rect 32 320 35 335
rect 22 315 26 316
rect 6 272 11 274
rect 6 2 8 272
rect 22 310 26 311
rect 22 305 26 306
rect 22 300 26 301
rect 22 295 26 296
rect 22 290 26 291
rect 22 285 26 286
rect 22 280 26 281
rect 30 319 35 320
rect 18 270 27 273
rect 34 316 35 319
rect 42 327 45 331
rect 53 327 56 346
rect 92 339 95 347
rect 98 347 115 348
rect 98 343 99 347
rect 107 343 108 347
rect 112 343 115 347
rect 98 342 115 343
rect 118 354 127 357
rect 135 364 139 365
rect 135 359 139 360
rect 139 355 151 357
rect 135 354 151 355
rect 64 331 83 332
rect 68 327 69 331
rect 73 327 74 331
rect 38 320 49 327
rect 64 323 83 327
rect 86 327 89 335
rect 98 331 115 332
rect 102 327 104 331
rect 108 327 109 331
rect 113 327 115 331
rect 98 326 115 327
rect 64 320 67 323
rect 78 321 83 323
rect 38 317 47 320
rect 46 316 47 317
rect 46 315 51 316
rect 46 311 47 315
rect 46 310 51 311
rect 46 306 47 310
rect 46 305 51 306
rect 46 301 47 305
rect 46 300 51 301
rect 46 296 47 300
rect 46 295 51 296
rect 46 291 47 295
rect 46 290 51 291
rect 46 286 47 290
rect 46 285 51 286
rect 46 281 47 285
rect 46 280 51 281
rect 46 276 47 280
rect 55 319 59 320
rect 43 270 55 273
rect 62 316 67 320
rect 62 312 63 316
rect 62 311 67 312
rect 62 307 63 311
rect 62 306 67 307
rect 62 302 63 306
rect 62 301 67 302
rect 62 297 63 301
rect 62 296 67 297
rect 62 292 63 296
rect 62 291 67 292
rect 62 287 63 291
rect 62 286 67 287
rect 62 282 63 286
rect 62 281 67 282
rect 62 277 63 281
rect 63 276 67 277
rect 59 270 60 274
rect 71 319 75 320
rect 24 267 27 270
rect 57 269 60 270
rect 78 317 79 321
rect 111 320 115 326
rect 78 316 83 317
rect 78 312 79 316
rect 78 311 83 312
rect 78 307 79 311
rect 78 306 83 307
rect 78 302 79 306
rect 78 301 83 302
rect 78 297 79 301
rect 78 296 83 297
rect 78 292 79 296
rect 78 291 83 292
rect 78 287 79 291
rect 78 286 83 287
rect 78 282 79 286
rect 78 281 83 282
rect 78 277 79 281
rect 78 276 83 277
rect 78 272 79 276
rect 71 269 75 270
rect 103 319 107 320
rect 94 316 99 318
rect 94 312 95 316
rect 94 311 99 312
rect 94 307 95 311
rect 94 306 99 307
rect 94 302 95 306
rect 94 301 99 302
rect 94 297 95 301
rect 94 296 99 297
rect 94 292 95 296
rect 94 291 99 292
rect 94 287 95 291
rect 94 286 99 287
rect 94 282 95 286
rect 94 281 99 282
rect 94 277 95 281
rect 94 276 99 277
rect 94 272 95 276
rect 87 269 91 271
rect 111 315 115 316
rect 118 320 121 354
rect 124 347 134 348
rect 128 343 130 347
rect 140 339 143 347
rect 127 327 130 335
rect 136 331 148 332
rect 136 327 137 331
rect 141 327 142 331
rect 146 327 148 331
rect 136 326 148 327
rect 151 320 154 353
rect 118 314 119 320
rect 111 310 115 311
rect 111 305 115 306
rect 111 300 115 301
rect 111 295 115 296
rect 111 290 115 291
rect 111 285 115 286
rect 111 280 115 281
rect 103 269 107 270
rect 110 271 119 273
rect 123 317 135 320
rect 135 314 139 316
rect 110 270 123 271
rect 127 311 131 313
rect 135 307 139 310
rect 131 272 143 275
rect 127 271 143 272
rect 147 317 154 320
rect 151 309 155 310
rect 110 269 114 270
rect 24 263 25 267
rect 57 266 114 269
rect 127 267 131 271
rect 117 264 131 267
rect 158 266 190 383
rect 218 380 221 383
rect 233 380 237 383
rect 249 383 285 386
rect 193 375 197 376
rect 193 370 197 371
rect 193 365 197 366
rect 193 360 197 361
rect 193 354 197 356
rect 205 377 217 380
rect 201 354 205 356
rect 209 364 213 365
rect 209 358 213 360
rect 194 348 197 354
rect 209 348 213 354
rect 194 346 213 348
rect 194 340 213 342
rect 217 354 221 356
rect 224 376 225 380
rect 224 375 229 376
rect 224 371 225 375
rect 224 370 229 371
rect 224 366 225 370
rect 224 365 229 366
rect 224 361 225 365
rect 224 360 229 361
rect 224 356 225 360
rect 224 354 229 356
rect 233 354 237 356
rect 241 380 245 382
rect 241 375 245 376
rect 241 370 245 371
rect 241 365 245 366
rect 241 360 245 361
rect 241 354 245 356
rect 249 380 253 383
rect 265 380 269 383
rect 281 380 285 383
rect 249 354 253 356
rect 257 375 261 376
rect 257 370 261 371
rect 257 365 261 366
rect 257 360 261 361
rect 217 339 220 354
rect 224 347 227 354
rect 242 348 245 354
rect 257 348 261 356
rect 194 331 213 332
rect 203 327 204 331
rect 208 327 209 331
rect 194 326 213 327
rect 194 318 197 326
rect 11 13 14 263
rect 17 258 36 260
rect 17 251 36 254
rect 17 240 36 243
rect 17 232 36 236
rect 26 228 36 232
rect 17 227 36 228
rect 26 226 36 227
rect 26 223 32 226
rect 17 222 32 223
rect 26 221 36 222
rect 39 242 42 257
rect 39 236 43 238
rect 26 208 29 221
rect 39 217 42 232
rect 17 207 29 208
rect 26 203 29 207
rect 17 202 29 203
rect 26 188 29 202
rect 17 187 29 188
rect 26 183 29 187
rect 17 182 29 183
rect 26 168 29 182
rect 17 167 29 168
rect 26 163 29 167
rect 17 162 29 163
rect 26 148 29 162
rect 17 147 29 148
rect 26 143 29 147
rect 17 142 29 143
rect 26 128 29 142
rect 17 127 29 128
rect 26 123 29 127
rect 17 122 29 123
rect 26 108 29 122
rect 17 107 29 108
rect 26 103 29 107
rect 17 102 29 103
rect 26 88 29 102
rect 17 87 29 88
rect 26 83 29 87
rect 17 82 29 83
rect 26 68 29 82
rect 17 67 29 68
rect 26 63 29 67
rect 17 62 29 63
rect 26 48 29 62
rect 17 47 29 48
rect 26 43 29 47
rect 36 214 42 217
rect 17 42 29 43
rect 26 37 29 42
rect 26 36 39 37
rect 26 33 32 36
rect 17 32 32 33
rect 36 33 39 36
rect 36 32 43 33
rect 17 31 43 32
rect 17 29 39 31
rect 21 25 23 29
rect 37 25 39 29
rect 17 24 39 25
rect 21 20 23 24
rect 37 23 39 24
rect 37 20 43 23
rect 17 19 43 20
rect 17 16 23 19
rect 37 16 43 19
rect 37 15 40 16
rect 23 14 40 15
rect 47 13 50 263
rect 57 260 59 263
rect 53 259 59 260
rect 113 259 114 263
rect 53 257 114 259
rect 53 253 54 257
rect 108 255 114 257
rect 53 251 107 253
rect 117 251 120 264
rect 134 261 190 266
rect 123 246 190 261
rect 193 316 197 318
rect 193 311 197 312
rect 193 306 197 307
rect 193 301 197 302
rect 193 291 197 292
rect 193 281 197 282
rect 193 276 197 277
rect 193 264 197 272
rect 201 316 205 320
rect 209 316 213 326
rect 209 311 213 312
rect 209 306 213 307
rect 209 301 213 302
rect 209 291 213 292
rect 209 281 213 282
rect 209 276 213 277
rect 217 320 220 335
rect 233 327 236 347
rect 242 346 261 348
rect 251 342 252 346
rect 256 342 257 346
rect 272 376 273 380
rect 272 375 277 376
rect 272 371 273 375
rect 272 370 277 371
rect 272 366 273 370
rect 272 365 277 366
rect 272 361 273 365
rect 272 360 277 361
rect 272 356 273 360
rect 242 331 261 332
rect 251 327 252 331
rect 256 327 257 331
rect 224 320 227 327
rect 242 326 261 327
rect 242 320 245 326
rect 217 316 221 320
rect 224 316 229 320
rect 224 312 225 316
rect 224 311 229 312
rect 224 307 225 311
rect 224 306 229 307
rect 224 302 225 306
rect 224 301 229 302
rect 224 292 225 301
rect 224 291 229 292
rect 224 282 225 291
rect 224 281 229 282
rect 224 277 225 281
rect 224 276 229 277
rect 224 272 225 276
rect 233 316 237 320
rect 201 267 205 272
rect 217 267 221 272
rect 233 267 237 272
rect 201 263 237 267
rect 193 258 230 260
rect 193 254 194 258
rect 228 254 230 258
rect 193 251 230 254
rect 193 247 194 251
rect 228 247 230 251
rect 233 250 237 263
rect 241 316 245 320
rect 241 311 245 312
rect 241 306 245 307
rect 241 301 245 302
rect 241 291 245 292
rect 241 281 245 282
rect 241 276 245 277
rect 241 265 245 272
rect 249 316 253 320
rect 257 316 261 326
rect 257 311 261 312
rect 257 306 261 307
rect 257 301 261 302
rect 257 291 261 292
rect 257 281 261 282
rect 257 276 261 277
rect 265 320 268 356
rect 272 355 277 356
rect 272 348 275 355
rect 281 354 285 356
rect 289 382 295 386
rect 299 382 300 386
rect 289 381 300 382
rect 289 380 295 381
rect 293 377 295 380
rect 299 377 300 381
rect 293 376 300 377
rect 289 375 295 376
rect 293 372 295 375
rect 299 372 300 376
rect 293 371 300 372
rect 289 370 295 371
rect 293 367 295 370
rect 299 367 300 371
rect 293 366 300 367
rect 289 365 295 366
rect 293 362 295 365
rect 299 362 300 366
rect 293 361 300 362
rect 289 360 295 361
rect 293 357 295 360
rect 299 357 300 361
rect 293 356 300 357
rect 289 354 295 356
rect 290 352 295 354
rect 299 352 300 356
rect 290 351 300 352
rect 271 346 275 348
rect 299 347 300 351
rect 280 339 283 347
rect 290 346 300 347
rect 299 342 300 346
rect 290 341 300 342
rect 271 331 275 332
rect 280 327 283 335
rect 271 326 275 327
rect 272 320 275 326
rect 290 323 295 332
rect 299 323 300 332
rect 290 321 300 323
rect 290 320 295 321
rect 265 316 269 320
rect 272 316 277 320
rect 272 312 273 316
rect 272 311 277 312
rect 272 307 273 311
rect 272 306 277 307
rect 272 302 273 306
rect 272 301 277 302
rect 272 292 273 301
rect 272 291 277 292
rect 272 282 273 291
rect 272 281 277 282
rect 272 277 273 281
rect 272 276 277 277
rect 272 272 273 276
rect 281 316 285 320
rect 249 267 253 272
rect 265 267 269 272
rect 281 267 285 272
rect 249 263 285 267
rect 289 316 295 320
rect 241 260 245 261
rect 240 259 254 260
rect 240 253 254 255
rect 233 246 253 250
rect 123 244 176 246
rect 53 241 120 243
rect 117 237 120 241
rect 53 233 120 237
rect 53 229 54 233
rect 63 229 64 233
rect 68 229 69 233
rect 78 229 79 233
rect 83 229 84 233
rect 93 229 94 233
rect 98 229 99 233
rect 108 229 109 233
rect 113 229 114 233
rect 118 229 120 233
rect 53 227 120 229
rect 53 223 54 227
rect 63 223 64 227
rect 68 223 69 227
rect 78 223 79 227
rect 83 223 84 227
rect 93 223 94 227
rect 98 223 99 227
rect 108 223 109 227
rect 113 223 114 227
rect 118 223 120 227
rect 53 214 120 223
rect 53 210 54 214
rect 118 210 120 214
rect 53 209 120 210
rect 123 205 143 244
rect 53 200 143 205
rect 53 196 56 200
rect 120 196 143 200
rect 53 194 143 196
rect 53 190 56 194
rect 120 190 143 194
rect 53 185 143 190
rect 53 181 120 182
rect 53 177 56 181
rect 53 167 120 177
rect 53 163 55 167
rect 64 163 65 167
rect 69 163 70 167
rect 79 163 80 167
rect 84 163 85 167
rect 94 163 95 167
rect 99 163 100 167
rect 109 163 110 167
rect 114 163 115 167
rect 119 163 120 167
rect 53 161 120 163
rect 53 157 55 161
rect 64 157 65 161
rect 69 157 70 161
rect 79 157 80 161
rect 84 157 85 161
rect 94 157 95 161
rect 99 157 100 161
rect 109 157 110 161
rect 114 157 115 161
rect 119 157 120 161
rect 53 148 120 157
rect 53 144 55 148
rect 119 144 120 148
rect 53 143 120 144
rect 123 139 143 185
rect 56 134 143 139
rect 120 125 143 134
rect 56 120 143 125
rect 53 116 120 117
rect 53 112 55 116
rect 119 112 120 116
rect 53 102 120 112
rect 53 98 54 102
rect 63 98 64 102
rect 68 98 69 102
rect 78 98 79 102
rect 83 98 84 102
rect 93 98 94 102
rect 98 98 99 102
rect 108 98 109 102
rect 113 98 114 102
rect 118 98 120 102
rect 53 96 120 98
rect 53 92 54 96
rect 63 92 64 96
rect 68 92 69 96
rect 78 92 79 96
rect 83 92 84 96
rect 93 92 94 96
rect 98 92 99 96
rect 108 92 109 96
rect 113 92 114 96
rect 118 92 120 96
rect 53 84 120 92
rect 53 80 55 84
rect 119 80 120 84
rect 53 78 120 80
rect 123 74 143 120
rect 53 69 143 74
rect 53 60 56 69
rect 120 60 143 69
rect 53 56 143 60
rect 53 51 119 52
rect 53 47 54 51
rect 118 47 119 51
rect 53 37 119 47
rect 57 33 59 37
rect 118 33 119 37
rect 53 32 119 33
rect 57 31 119 32
rect 57 17 59 31
rect 63 17 64 31
rect 68 17 69 31
rect 73 17 74 31
rect 78 17 79 31
rect 83 17 84 31
rect 88 17 89 31
rect 93 17 94 31
rect 98 17 99 31
rect 103 17 104 31
rect 108 17 109 31
rect 113 17 114 31
rect 118 17 119 31
rect 57 14 119 17
rect 123 49 143 56
rect 147 239 153 240
rect 147 230 148 239
rect 152 230 153 239
rect 147 229 153 230
rect 147 225 148 229
rect 152 225 153 229
rect 147 224 153 225
rect 147 215 148 224
rect 152 215 153 224
rect 147 214 153 215
rect 147 210 148 214
rect 152 210 153 214
rect 147 209 153 210
rect 147 200 148 209
rect 152 200 153 209
rect 147 199 153 200
rect 147 195 148 199
rect 152 195 153 199
rect 147 194 153 195
rect 147 185 148 194
rect 152 185 153 194
rect 147 184 153 185
rect 147 180 148 184
rect 152 180 153 184
rect 147 179 153 180
rect 147 170 148 179
rect 152 170 153 179
rect 147 169 153 170
rect 147 165 148 169
rect 152 165 153 169
rect 147 164 153 165
rect 147 155 148 164
rect 152 155 153 164
rect 147 154 153 155
rect 147 150 148 154
rect 152 150 153 154
rect 147 144 153 150
rect 147 140 148 144
rect 152 140 153 144
rect 147 139 153 140
rect 147 135 148 139
rect 152 135 153 139
rect 147 134 153 135
rect 147 125 148 134
rect 152 125 153 134
rect 147 124 153 125
rect 147 120 148 124
rect 152 120 153 124
rect 147 119 153 120
rect 147 110 148 119
rect 152 110 153 119
rect 147 109 153 110
rect 147 105 148 109
rect 152 105 153 109
rect 147 104 153 105
rect 147 95 148 104
rect 152 95 153 104
rect 147 94 153 95
rect 147 90 148 94
rect 152 90 153 94
rect 147 89 153 90
rect 147 85 148 89
rect 152 85 153 89
rect 147 79 153 85
rect 147 75 148 79
rect 152 75 153 79
rect 147 74 153 75
rect 147 65 148 74
rect 152 65 153 74
rect 147 64 153 65
rect 147 60 148 64
rect 152 60 153 64
rect 147 59 153 60
rect 147 55 148 59
rect 152 55 153 59
rect 147 54 153 55
rect 157 205 176 244
rect 179 241 247 243
rect 179 237 182 241
rect 246 237 247 241
rect 179 233 247 237
rect 179 229 182 233
rect 191 229 192 233
rect 196 229 197 233
rect 206 229 207 233
rect 211 229 212 233
rect 221 229 222 233
rect 226 229 227 233
rect 236 229 237 233
rect 241 229 242 233
rect 246 229 247 233
rect 179 227 247 229
rect 179 223 182 227
rect 191 223 192 227
rect 196 223 197 227
rect 206 223 207 227
rect 211 223 212 227
rect 221 223 222 227
rect 226 223 227 227
rect 236 223 237 227
rect 241 223 242 227
rect 246 223 247 227
rect 179 214 247 223
rect 179 210 182 214
rect 246 210 247 214
rect 179 209 247 210
rect 157 200 247 205
rect 157 196 180 200
rect 244 196 247 200
rect 157 194 247 196
rect 157 190 180 194
rect 244 190 247 194
rect 157 185 247 190
rect 157 139 176 185
rect 180 181 247 182
rect 180 177 182 181
rect 246 177 247 181
rect 180 167 247 177
rect 180 163 181 167
rect 190 163 191 167
rect 195 163 196 167
rect 205 163 206 167
rect 210 163 211 167
rect 220 163 221 167
rect 225 163 226 167
rect 235 163 236 167
rect 240 163 241 167
rect 245 163 247 167
rect 180 161 247 163
rect 180 157 181 161
rect 190 157 191 161
rect 195 157 196 161
rect 205 157 206 161
rect 210 157 211 161
rect 220 157 221 161
rect 225 157 226 161
rect 235 157 236 161
rect 240 157 241 161
rect 245 157 247 161
rect 180 148 247 157
rect 180 144 181 148
rect 245 144 247 148
rect 180 143 247 144
rect 157 134 247 139
rect 157 125 180 134
rect 244 125 247 134
rect 157 120 247 125
rect 157 74 176 120
rect 180 115 247 117
rect 180 111 182 115
rect 246 111 247 115
rect 180 102 247 111
rect 180 98 182 102
rect 191 98 192 102
rect 196 98 197 102
rect 206 98 207 102
rect 211 98 212 102
rect 221 98 222 102
rect 226 98 227 102
rect 236 98 237 102
rect 241 98 242 102
rect 246 98 247 102
rect 180 96 247 98
rect 180 92 182 96
rect 191 92 192 96
rect 196 92 197 96
rect 206 92 207 96
rect 211 92 212 96
rect 221 92 222 96
rect 226 92 227 96
rect 236 92 237 96
rect 241 92 242 96
rect 246 92 247 96
rect 180 84 247 92
rect 180 80 182 84
rect 246 80 247 84
rect 180 78 247 80
rect 157 69 247 74
rect 157 60 180 69
rect 244 60 247 69
rect 157 56 247 60
rect 157 49 176 56
rect 123 19 176 49
rect 123 15 128 19
rect 172 15 176 19
rect 123 12 176 15
rect 180 51 247 52
rect 180 47 182 51
rect 246 47 247 51
rect 180 37 247 47
rect 180 33 182 37
rect 246 33 247 37
rect 180 31 247 33
rect 180 17 182 31
rect 186 17 187 31
rect 191 17 192 31
rect 196 17 197 31
rect 201 17 202 31
rect 206 17 207 31
rect 211 17 212 31
rect 216 17 217 31
rect 221 17 222 31
rect 226 17 227 31
rect 231 17 232 31
rect 236 17 237 31
rect 241 17 242 31
rect 246 17 247 31
rect 180 16 247 17
rect 180 14 241 16
rect 250 13 253 246
rect 257 13 260 263
rect 287 257 289 260
rect 293 257 295 316
rect 299 257 300 321
rect 287 256 300 257
rect 263 251 300 256
rect 287 247 290 251
rect 263 236 267 238
rect 264 217 267 232
rect 274 229 276 243
rect 271 228 276 229
rect 263 36 271 37
rect 263 32 264 36
rect 268 32 271 36
rect 263 30 271 32
rect 267 16 271 30
rect 269 14 271 16
rect 275 14 276 228
rect 280 228 286 243
rect 280 14 282 228
rect 289 8 290 247
rect 56 6 241 8
rect 269 6 290 8
rect 287 2 290 6
rect 299 2 300 251
rect 0 0 300 2
<< m2contact >>
rect 14 440 18 654
rect 22 650 111 654
rect 22 641 26 645
rect 30 631 44 645
rect 61 631 65 645
rect 76 631 80 645
rect 91 631 95 645
rect 106 631 110 645
rect 20 621 29 625
rect 32 621 36 625
rect 20 601 29 605
rect 20 581 29 585
rect 20 561 29 565
rect 32 555 36 589
rect 41 587 50 621
rect 52 618 116 622
rect 52 586 116 590
rect 41 572 60 576
rect 71 572 75 576
rect 86 572 90 576
rect 101 572 105 576
rect 41 566 60 570
rect 71 566 75 570
rect 86 566 90 570
rect 101 566 105 570
rect 20 541 29 545
rect 20 521 29 525
rect 20 501 29 505
rect 32 490 36 524
rect 42 522 51 556
rect 55 552 114 556
rect 55 522 114 526
rect 41 508 60 512
rect 71 508 75 512
rect 86 508 90 512
rect 101 508 105 512
rect 41 502 60 506
rect 71 502 75 506
rect 86 502 90 506
rect 101 502 105 506
rect 20 481 29 485
rect 20 461 29 465
rect 20 441 29 445
rect 42 458 51 492
rect 55 489 114 493
rect 54 457 113 461
rect 40 443 49 447
rect 51 443 60 447
rect 71 443 75 447
rect 86 443 90 447
rect 101 443 105 447
rect 46 437 50 441
rect 56 437 60 441
rect 71 437 75 441
rect 86 437 90 441
rect 101 437 105 441
rect 32 431 41 435
rect 15 421 29 425
rect 7 395 11 409
rect 13 405 27 409
rect 39 421 113 425
rect 39 405 108 409
rect 148 638 152 642
rect 148 618 152 622
rect 148 598 152 602
rect 148 578 152 582
rect 148 558 152 562
rect 148 538 152 542
rect 148 518 152 522
rect 148 498 152 502
rect 148 478 152 482
rect 148 458 152 462
rect 148 438 152 442
rect 189 651 278 655
rect 188 631 192 645
rect 203 631 207 645
rect 218 631 222 645
rect 233 631 237 645
rect 254 631 268 645
rect 271 641 280 645
rect 186 618 245 622
rect 264 621 268 625
rect 271 621 280 625
rect 186 585 245 589
rect 249 586 258 620
rect 271 601 280 605
rect 194 572 198 576
rect 209 572 213 576
rect 224 572 228 576
rect 239 572 258 576
rect 194 566 198 570
rect 209 566 213 570
rect 224 566 228 570
rect 239 566 258 570
rect 186 553 245 557
rect 186 522 245 526
rect 249 522 258 556
rect 264 554 268 588
rect 271 581 280 585
rect 271 561 280 565
rect 271 541 280 545
rect 193 508 197 512
rect 208 508 212 512
rect 223 508 227 512
rect 238 508 257 512
rect 193 502 197 506
rect 208 502 212 506
rect 223 502 227 506
rect 238 502 257 506
rect 184 489 248 493
rect 148 421 152 425
rect 187 457 246 461
rect 250 458 259 492
rect 264 490 268 524
rect 271 521 280 525
rect 271 501 280 505
rect 194 443 198 447
rect 209 443 213 447
rect 224 443 228 447
rect 239 443 243 447
rect 245 443 254 447
rect 256 443 260 447
rect 194 437 198 441
rect 209 437 213 441
rect 224 437 228 441
rect 239 437 243 441
rect 249 437 253 441
rect 259 431 268 435
rect 271 481 280 485
rect 271 461 280 465
rect 271 441 280 445
rect 282 441 286 655
rect 184 421 288 425
rect 295 407 299 411
rect 7 354 11 393
rect 295 397 299 401
rect 289 388 293 392
rect 295 387 299 391
rect 22 371 26 375
rect 22 361 26 365
rect 47 369 51 373
rect 47 359 51 363
rect 63 369 67 373
rect 63 359 67 363
rect 79 369 83 373
rect 79 359 83 363
rect 95 369 99 373
rect 95 359 99 363
rect 111 369 115 373
rect 111 359 115 363
rect 119 360 123 364
rect 20 335 29 339
rect 7 274 11 318
rect 22 311 26 315
rect 22 301 26 305
rect 22 291 26 295
rect 22 281 26 285
rect 103 343 107 347
rect 135 360 139 364
rect 92 335 101 339
rect 69 327 73 331
rect 104 327 108 331
rect 47 311 51 315
rect 47 301 51 305
rect 47 291 51 295
rect 47 281 51 285
rect 63 307 67 311
rect 63 297 67 301
rect 63 287 67 291
rect 63 277 67 281
rect 79 317 83 321
rect 79 307 83 311
rect 79 297 83 301
rect 79 287 83 291
rect 79 277 83 281
rect 95 307 99 311
rect 95 297 99 301
rect 95 287 99 291
rect 95 277 99 281
rect 111 311 115 315
rect 130 343 134 347
rect 124 335 133 339
rect 142 327 146 331
rect 111 301 115 305
rect 111 291 115 295
rect 111 281 115 285
rect 135 310 139 314
rect 151 310 155 314
rect 193 371 197 375
rect 193 361 197 365
rect 209 360 213 364
rect 194 336 213 340
rect 225 371 229 375
rect 225 361 229 365
rect 241 371 245 375
rect 241 361 245 365
rect 257 371 261 375
rect 257 361 261 365
rect 217 335 226 339
rect 204 327 208 331
rect 17 247 36 251
rect 17 223 26 227
rect 32 222 36 226
rect 39 238 43 242
rect 39 232 43 236
rect 17 203 26 207
rect 17 183 26 187
rect 17 163 26 167
rect 17 143 26 147
rect 17 123 26 127
rect 17 103 26 107
rect 17 83 26 87
rect 17 63 26 67
rect 17 43 26 47
rect 32 32 36 36
rect 17 20 21 24
rect 23 20 37 24
rect 39 23 43 27
rect 53 247 107 251
rect 111 247 120 251
rect 193 307 197 311
rect 193 292 197 301
rect 193 277 197 281
rect 209 307 213 311
rect 209 292 213 301
rect 209 277 213 281
rect 252 342 256 346
rect 273 371 277 375
rect 273 361 277 365
rect 252 327 256 331
rect 225 307 229 311
rect 225 292 229 301
rect 225 277 229 281
rect 194 247 228 251
rect 241 307 245 311
rect 241 292 245 301
rect 241 277 245 281
rect 257 307 261 311
rect 257 292 261 301
rect 257 277 261 281
rect 295 377 299 381
rect 289 371 293 375
rect 295 367 299 371
rect 289 361 293 365
rect 295 357 299 361
rect 290 347 299 351
rect 277 335 286 339
rect 273 307 277 311
rect 273 292 277 301
rect 273 277 277 281
rect 64 229 68 233
rect 79 229 83 233
rect 94 229 98 233
rect 109 229 113 233
rect 64 223 68 227
rect 79 223 83 227
rect 94 223 98 227
rect 109 223 113 227
rect 54 210 118 214
rect 56 177 120 181
rect 65 163 69 167
rect 80 163 84 167
rect 95 163 99 167
rect 110 163 114 167
rect 65 157 69 161
rect 80 157 84 161
rect 95 157 99 161
rect 110 157 114 161
rect 55 144 119 148
rect 55 112 119 116
rect 64 98 68 102
rect 79 98 83 102
rect 94 98 98 102
rect 109 98 113 102
rect 64 92 68 96
rect 79 92 83 96
rect 94 92 98 96
rect 109 92 113 96
rect 55 80 119 84
rect 54 47 118 51
rect 59 17 63 31
rect 69 17 73 31
rect 79 17 83 31
rect 89 17 93 31
rect 99 17 103 31
rect 109 17 113 31
rect 148 225 152 229
rect 148 210 152 214
rect 148 195 152 199
rect 148 180 152 184
rect 148 165 152 169
rect 148 150 152 154
rect 148 135 152 139
rect 148 120 152 124
rect 148 105 152 109
rect 148 90 152 94
rect 148 75 152 79
rect 148 60 152 64
rect 192 229 196 233
rect 207 229 211 233
rect 222 229 226 233
rect 237 229 241 233
rect 192 223 196 227
rect 207 223 211 227
rect 222 223 226 227
rect 237 223 241 227
rect 182 210 246 214
rect 182 177 246 181
rect 191 163 195 167
rect 206 163 210 167
rect 221 163 225 167
rect 236 163 240 167
rect 191 157 195 161
rect 206 157 210 161
rect 221 157 225 161
rect 236 157 240 161
rect 181 144 245 148
rect 182 111 246 115
rect 192 98 196 102
rect 207 98 211 102
rect 222 98 226 102
rect 237 98 241 102
rect 192 92 196 96
rect 207 92 211 96
rect 222 92 226 96
rect 237 92 241 96
rect 182 80 246 84
rect 128 15 172 19
rect 11 9 20 13
rect 44 9 53 13
rect 182 47 246 51
rect 187 17 191 31
rect 197 17 201 31
rect 207 17 211 31
rect 217 17 221 31
rect 227 17 231 31
rect 237 17 241 31
rect 244 9 253 13
rect 295 257 299 321
rect 263 247 287 251
rect 263 238 267 242
rect 263 232 267 236
rect 264 32 268 36
rect 271 14 275 228
rect 282 14 286 228
rect 257 9 266 13
<< metal2 >>
rect 20 997 280 1000
rect 20 743 23 997
rect 277 743 280 997
rect 20 740 280 743
rect 0 655 300 670
rect 0 654 189 655
rect 0 440 14 654
rect 18 650 22 654
rect 111 651 189 654
rect 278 651 282 655
rect 111 650 282 651
rect 18 645 282 650
rect 18 641 22 645
rect 26 641 30 645
rect 18 631 30 641
rect 44 631 61 645
rect 65 631 76 645
rect 80 631 91 645
rect 95 631 106 645
rect 110 642 188 645
rect 110 638 148 642
rect 152 638 188 642
rect 110 631 188 638
rect 192 631 203 645
rect 207 631 218 645
rect 222 631 233 645
rect 237 631 254 645
rect 268 641 271 645
rect 280 641 282 645
rect 268 631 282 641
rect 18 625 282 631
rect 18 621 20 625
rect 29 621 32 625
rect 36 622 264 625
rect 36 621 52 622
rect 18 605 41 621
rect 18 601 20 605
rect 29 601 41 605
rect 18 589 41 601
rect 18 585 32 589
rect 18 581 20 585
rect 29 581 32 585
rect 18 565 32 581
rect 18 561 20 565
rect 29 561 32 565
rect 18 555 32 561
rect 36 587 41 589
rect 50 618 52 621
rect 116 618 148 622
rect 152 618 186 622
rect 245 621 264 622
rect 268 621 271 625
rect 280 621 282 625
rect 245 620 282 621
rect 245 618 249 620
rect 50 602 249 618
rect 50 598 148 602
rect 152 598 249 602
rect 50 590 249 598
rect 50 587 52 590
rect 36 586 52 587
rect 116 589 249 590
rect 116 586 186 589
rect 36 585 186 586
rect 245 586 249 589
rect 258 605 282 620
rect 258 601 271 605
rect 280 601 282 605
rect 258 588 282 601
rect 258 586 264 588
rect 245 585 264 586
rect 36 582 264 585
rect 36 578 148 582
rect 152 578 264 582
rect 36 576 264 578
rect 36 572 41 576
rect 60 572 71 576
rect 75 572 86 576
rect 90 572 101 576
rect 105 572 194 576
rect 198 572 209 576
rect 213 572 224 576
rect 228 572 239 576
rect 258 572 264 576
rect 36 570 264 572
rect 36 566 41 570
rect 60 566 71 570
rect 75 566 86 570
rect 90 566 101 570
rect 105 566 194 570
rect 198 566 209 570
rect 213 566 224 570
rect 228 566 239 570
rect 258 566 264 570
rect 36 562 264 566
rect 36 558 148 562
rect 152 558 264 562
rect 36 557 264 558
rect 36 556 186 557
rect 36 555 42 556
rect 18 545 42 555
rect 18 541 20 545
rect 29 541 42 545
rect 18 525 42 541
rect 18 521 20 525
rect 29 524 42 525
rect 29 521 32 524
rect 18 505 32 521
rect 18 501 20 505
rect 29 501 32 505
rect 18 490 32 501
rect 36 522 42 524
rect 51 552 55 556
rect 114 553 186 556
rect 245 556 264 557
rect 245 553 249 556
rect 114 552 249 553
rect 51 542 249 552
rect 51 538 148 542
rect 152 538 249 542
rect 51 526 249 538
rect 51 522 55 526
rect 114 522 186 526
rect 245 522 249 526
rect 258 554 264 556
rect 268 585 282 588
rect 268 581 271 585
rect 280 581 282 585
rect 268 565 282 581
rect 268 561 271 565
rect 280 561 282 565
rect 268 554 282 561
rect 258 545 282 554
rect 258 541 271 545
rect 280 541 282 545
rect 258 525 282 541
rect 258 524 271 525
rect 258 522 264 524
rect 36 518 148 522
rect 152 518 264 522
rect 36 512 264 518
rect 36 508 41 512
rect 60 508 71 512
rect 75 508 86 512
rect 90 508 101 512
rect 105 508 193 512
rect 197 508 208 512
rect 212 508 223 512
rect 227 508 238 512
rect 257 508 264 512
rect 36 506 264 508
rect 36 502 41 506
rect 60 502 71 506
rect 75 502 86 506
rect 90 502 101 506
rect 105 502 193 506
rect 197 502 208 506
rect 212 502 223 506
rect 227 502 238 506
rect 257 502 264 506
rect 36 498 148 502
rect 152 498 264 502
rect 36 493 264 498
rect 36 492 55 493
rect 36 490 42 492
rect 18 485 42 490
rect 18 481 20 485
rect 29 481 42 485
rect 18 465 42 481
rect 18 461 20 465
rect 29 461 42 465
rect 18 458 42 461
rect 51 489 55 492
rect 114 489 184 493
rect 248 492 264 493
rect 248 489 250 492
rect 51 482 250 489
rect 51 478 148 482
rect 152 478 250 482
rect 51 462 250 478
rect 51 461 148 462
rect 51 458 54 461
rect 18 457 54 458
rect 113 458 148 461
rect 152 461 250 462
rect 152 458 187 461
rect 113 457 187 458
rect 246 458 250 461
rect 259 490 264 492
rect 268 521 271 524
rect 280 521 282 525
rect 268 505 282 521
rect 268 501 271 505
rect 280 501 282 505
rect 268 490 282 501
rect 259 485 282 490
rect 259 481 271 485
rect 280 481 282 485
rect 259 465 282 481
rect 259 461 271 465
rect 280 461 282 465
rect 259 458 282 461
rect 246 457 282 458
rect 18 447 282 457
rect 18 445 40 447
rect 18 441 20 445
rect 29 443 40 445
rect 49 443 51 447
rect 60 443 71 447
rect 75 443 86 447
rect 90 443 101 447
rect 105 443 194 447
rect 198 443 209 447
rect 213 443 224 447
rect 228 443 239 447
rect 243 443 245 447
rect 254 443 256 447
rect 260 445 282 447
rect 260 443 271 445
rect 29 442 271 443
rect 29 441 148 442
rect 18 440 46 441
rect 0 439 29 440
rect 45 437 46 440
rect 50 437 56 441
rect 60 437 71 441
rect 75 437 86 441
rect 90 437 101 441
rect 105 438 148 441
rect 152 441 271 442
rect 280 441 282 445
rect 286 441 300 655
rect 152 438 194 441
rect 105 437 194 438
rect 198 437 209 441
rect 213 437 224 441
rect 228 437 239 441
rect 243 437 249 441
rect 253 440 300 441
rect 253 437 255 440
rect 271 439 300 440
rect 32 435 41 436
rect 259 435 268 436
rect 41 431 259 433
rect 32 430 268 431
rect 36 429 268 430
rect 10 422 15 425
rect 0 421 15 422
rect 29 421 39 425
rect 113 421 148 425
rect 152 421 184 425
rect 288 421 300 422
rect 0 411 300 421
rect 0 409 295 411
rect 0 395 7 409
rect 11 405 13 409
rect 27 405 39 409
rect 108 407 295 409
rect 299 407 300 411
rect 108 405 300 407
rect 11 401 300 405
rect 11 397 295 401
rect 299 397 300 401
rect 11 395 300 397
rect 0 393 300 395
rect 0 354 7 393
rect 11 392 300 393
rect 11 388 289 392
rect 293 391 300 392
rect 293 388 295 391
rect 11 387 295 388
rect 299 387 300 391
rect 11 381 300 387
rect 11 377 295 381
rect 299 377 300 381
rect 11 375 300 377
rect 11 371 22 375
rect 26 373 193 375
rect 26 371 47 373
rect 11 369 47 371
rect 51 369 63 373
rect 67 369 79 373
rect 83 369 95 373
rect 99 369 111 373
rect 115 371 193 373
rect 197 371 225 375
rect 229 371 241 375
rect 245 371 257 375
rect 261 371 273 375
rect 277 371 289 375
rect 293 371 300 375
rect 115 369 295 371
rect 11 368 295 369
rect 11 365 115 368
rect 11 361 22 365
rect 26 363 115 365
rect 143 367 295 368
rect 299 367 300 371
rect 143 365 300 367
rect 26 361 47 363
rect 11 359 47 361
rect 51 359 63 363
rect 67 359 79 363
rect 83 359 95 363
rect 99 359 111 363
rect 123 360 135 364
rect 143 361 193 365
rect 197 364 225 365
rect 197 361 209 364
rect 143 360 209 361
rect 213 361 225 364
rect 229 361 241 365
rect 245 361 257 365
rect 261 361 273 365
rect 277 361 289 365
rect 293 361 300 365
rect 213 360 295 361
rect 11 355 115 359
rect 143 357 295 360
rect 299 357 300 361
rect 143 355 300 357
rect 11 354 300 355
rect 0 351 300 354
rect 0 347 290 351
rect 299 347 300 351
rect 0 343 103 347
rect 107 343 130 347
rect 134 346 300 347
rect 134 343 252 346
rect 136 341 213 343
rect 242 342 252 343
rect 256 343 300 346
rect 256 342 261 343
rect 194 340 213 341
rect 29 335 92 338
rect 101 335 124 338
rect 226 335 277 338
rect 136 331 213 332
rect 8 327 69 331
rect 73 327 104 331
rect 108 327 115 331
rect 8 326 115 327
rect 136 327 142 331
rect 146 327 204 331
rect 208 329 213 331
rect 242 329 252 331
rect 208 327 252 329
rect 256 327 261 331
rect 136 326 261 327
rect 0 321 300 326
rect 0 318 79 321
rect 0 274 7 318
rect 11 317 79 318
rect 83 318 295 321
rect 83 317 131 318
rect 11 315 131 317
rect 11 311 22 315
rect 26 311 47 315
rect 51 311 111 315
rect 115 311 131 315
rect 11 307 63 311
rect 67 307 79 311
rect 83 307 95 311
rect 99 307 131 311
rect 139 310 151 314
rect 159 311 295 318
rect 11 306 131 307
rect 159 307 193 311
rect 197 307 209 311
rect 213 307 225 311
rect 229 307 241 311
rect 245 307 257 311
rect 261 307 273 311
rect 277 307 295 311
rect 159 306 295 307
rect 11 305 295 306
rect 11 301 22 305
rect 26 301 47 305
rect 51 301 111 305
rect 115 301 295 305
rect 11 297 63 301
rect 67 297 79 301
rect 83 297 95 301
rect 99 297 193 301
rect 11 295 193 297
rect 11 291 22 295
rect 26 291 47 295
rect 51 291 111 295
rect 115 292 193 295
rect 197 292 209 301
rect 213 292 225 301
rect 229 292 241 301
rect 245 292 257 301
rect 261 292 273 301
rect 277 292 295 301
rect 115 291 295 292
rect 11 287 63 291
rect 67 287 79 291
rect 83 287 95 291
rect 99 287 295 291
rect 11 285 295 287
rect 11 281 22 285
rect 26 281 47 285
rect 51 281 111 285
rect 115 281 295 285
rect 11 277 63 281
rect 67 277 79 281
rect 83 277 95 281
rect 99 277 193 281
rect 197 277 209 281
rect 213 277 225 281
rect 229 277 241 281
rect 245 277 257 281
rect 261 277 273 281
rect 277 277 295 281
rect 11 274 295 277
rect 0 257 295 274
rect 299 257 300 321
rect 0 255 300 257
rect 0 253 108 255
rect 0 251 107 253
rect 124 251 300 255
rect 0 247 17 251
rect 36 247 53 251
rect 0 246 107 247
rect 111 242 120 247
rect 124 247 194 251
rect 228 247 263 251
rect 287 247 300 251
rect 124 246 300 247
rect 43 238 263 242
rect 39 236 43 238
rect 263 236 267 238
rect 0 228 35 230
rect 54 229 64 233
rect 68 229 79 233
rect 83 229 94 233
rect 98 229 109 233
rect 113 229 192 233
rect 196 229 207 233
rect 211 229 222 233
rect 226 229 237 233
rect 241 229 246 233
rect 54 228 148 229
rect 0 227 148 228
rect 0 223 17 227
rect 26 226 64 227
rect 26 223 32 226
rect 0 222 32 223
rect 36 223 64 226
rect 68 223 79 227
rect 83 223 94 227
rect 98 223 109 227
rect 113 225 148 227
rect 152 228 246 229
rect 280 228 300 230
rect 152 227 271 228
rect 152 225 192 227
rect 113 223 192 225
rect 196 223 207 227
rect 211 223 222 227
rect 226 223 237 227
rect 241 223 271 227
rect 36 222 271 223
rect 0 214 271 222
rect 0 210 54 214
rect 118 210 148 214
rect 152 210 182 214
rect 246 210 271 214
rect 0 207 271 210
rect 0 203 17 207
rect 26 203 271 207
rect 0 199 271 203
rect 0 195 148 199
rect 152 195 271 199
rect 0 187 271 195
rect 0 183 17 187
rect 26 184 271 187
rect 26 183 148 184
rect 0 181 148 183
rect 0 177 56 181
rect 120 180 148 181
rect 152 181 271 184
rect 152 180 182 181
rect 120 177 182 180
rect 246 177 271 181
rect 0 169 271 177
rect 0 167 148 169
rect 0 163 17 167
rect 26 163 65 167
rect 69 163 80 167
rect 84 163 95 167
rect 99 163 110 167
rect 114 165 148 167
rect 152 167 271 169
rect 152 165 191 167
rect 114 163 191 165
rect 195 163 206 167
rect 210 163 221 167
rect 225 163 236 167
rect 240 163 271 167
rect 0 161 271 163
rect 0 157 65 161
rect 69 157 80 161
rect 84 157 95 161
rect 99 157 110 161
rect 114 157 191 161
rect 195 157 206 161
rect 210 157 221 161
rect 225 157 236 161
rect 240 157 271 161
rect 0 154 271 157
rect 0 150 148 154
rect 152 150 271 154
rect 0 148 271 150
rect 0 147 55 148
rect 0 143 17 147
rect 26 144 55 147
rect 119 144 181 148
rect 245 144 271 148
rect 26 143 271 144
rect 0 139 271 143
rect 0 135 148 139
rect 152 135 271 139
rect 0 127 271 135
rect 0 123 17 127
rect 26 124 271 127
rect 26 123 148 124
rect 0 120 148 123
rect 152 120 271 124
rect 0 116 271 120
rect 0 112 55 116
rect 119 115 271 116
rect 119 112 182 115
rect 0 111 182 112
rect 246 111 271 115
rect 0 109 271 111
rect 0 107 148 109
rect 0 103 17 107
rect 26 105 148 107
rect 152 105 271 109
rect 26 103 271 105
rect 0 102 271 103
rect 0 98 64 102
rect 68 98 79 102
rect 83 98 94 102
rect 98 98 109 102
rect 113 98 192 102
rect 196 98 207 102
rect 211 98 222 102
rect 226 98 237 102
rect 241 98 271 102
rect 0 96 271 98
rect 0 92 64 96
rect 68 92 79 96
rect 83 92 94 96
rect 98 92 109 96
rect 113 94 192 96
rect 113 92 148 94
rect 0 90 148 92
rect 152 92 192 94
rect 196 92 207 96
rect 211 92 222 96
rect 226 92 237 96
rect 241 92 271 96
rect 152 90 271 92
rect 0 87 271 90
rect 0 83 17 87
rect 26 84 271 87
rect 26 83 55 84
rect 0 80 55 83
rect 119 80 182 84
rect 246 80 271 84
rect 0 79 271 80
rect 0 75 148 79
rect 152 75 271 79
rect 0 67 271 75
rect 0 63 17 67
rect 26 64 271 67
rect 26 63 148 64
rect 0 60 148 63
rect 152 60 271 64
rect 0 51 271 60
rect 0 47 54 51
rect 118 47 182 51
rect 246 47 271 51
rect 0 43 17 47
rect 26 43 271 47
rect 0 36 271 43
rect 0 32 32 36
rect 36 32 264 36
rect 268 32 271 36
rect 0 31 271 32
rect 0 27 59 31
rect 0 24 39 27
rect 0 20 17 24
rect 21 20 23 24
rect 37 23 39 24
rect 43 23 59 27
rect 37 20 59 23
rect 0 19 59 20
rect 0 0 7 19
rect 23 15 40 19
rect 11 0 20 9
rect 24 0 40 15
rect 57 17 59 19
rect 63 17 69 31
rect 73 17 79 31
rect 83 17 89 31
rect 93 17 99 31
rect 103 17 109 31
rect 113 23 187 31
rect 113 17 123 23
rect 44 0 53 9
rect 57 0 123 17
rect 128 0 172 15
rect 176 17 187 23
rect 191 17 197 31
rect 201 17 207 31
rect 211 17 217 31
rect 221 17 227 31
rect 231 17 237 31
rect 241 17 271 31
rect 176 0 240 17
rect 263 16 267 17
rect 270 14 271 17
rect 275 14 282 228
rect 286 14 300 228
rect 244 0 253 9
rect 257 0 266 9
rect 270 0 300 14
<< pad >>
rect 23 743 277 997
<< pseudo_rpoly >>
rect 126 405 191 407
rect 210 405 274 407
rect 126 393 191 395
rect 210 393 274 395
<< rpoly >>
rect 126 395 191 405
rect 210 395 274 405
<< m2p >>
rect 13 -2 17 2
rect 46 -2 50 2
rect 259 -2 263 2
<< m3p >>
rect 127 842 145 859
<< labels >>
rlabel metal2 48 0 48 0 8 DO
rlabel metal2 261 0 261 0 8 DI
rlabel metal2 15 0 15 0 1 OEN
rlabel metal2 169 129 169 129 1 Gnd2
rlabel metal2 132 535 132 535 1 Vdd2
rlabel metal2 174 307 174 307 1 Vdd
rlabel metal2 171 364 171 364 1 Gnd
rlabel m3p 136 850 136 850 1 YPAD
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1697747334
<< locali >>
rect 2 476 11 545
rect 232 476 268 546
rect 198 301 199 302
rect 2 226 76 301
rect 198 226 296 301
rect 416 226 508 290
rect 218 -8 256 60
rect 499 -8 508 61
use inv  inv_0
timestamp 1695393163
transform 1 0 124 0 1 151
box -122 -159 166 448
use inv  inv_1
timestamp 1695393163
transform 1 0 342 0 1 151
box -122 -159 166 448
<< labels >>
rlabel locali 26 262 26 262 0 A
port 1 e
rlabel locali 460 260 460 260 0 Y
port 2 w
rlabel locali 244 512 244 512 0 vdd
port 3 n
rlabel locali 236 26 236 26 1 gnd
port 4 n
<< end >>

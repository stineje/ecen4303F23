magic
tech scmos
magscale 1 30
timestamp 1160594422
<< error_p >>
rect 5130 44250 5760 44310
rect 11280 44250 12480 44310
rect 12720 44250 13920 44310
rect 14400 44250 15600 44310
rect 15750 44250 17280 44310
rect 17760 44250 19440 44310
rect 21360 44250 22800 44310
rect 24000 44250 25200 44310
rect 25680 44250 26880 44310
rect 27030 44250 28080 44310
rect 29430 44250 30480 44310
rect 30960 44250 31920 44310
rect 32400 44250 33450 44310
rect 33600 44250 34800 44310
rect 35040 44250 36000 44310
rect 38400 44250 39600 44310
rect 40800 44250 43200 44310
rect 48720 44250 50310 44310
rect 5130 38250 5730 38310
rect 6840 38250 8130 38310
rect 9000 38250 9480 38310
rect 20280 38250 20850 38310
rect 25800 38250 26100 38310
rect 27480 38250 27720 38310
rect 28440 38250 29280 38310
rect 37080 38250 37650 38310
rect 38520 38250 38760 38310
rect 39960 38250 40080 38310
rect 41070 38250 41640 38310
rect 44040 38250 44520 38310
rect 45240 38250 45720 38310
rect 46920 38250 47400 38310
rect 48600 38250 49170 38310
rect 50040 38250 50310 38310
rect 5130 32250 5520 32310
rect 10680 32250 10920 32310
rect 12840 32250 13560 32310
rect 14280 32250 14880 32310
rect 16080 32250 16440 32310
rect 18480 32250 19170 32310
rect 22800 32250 23160 32310
rect 24360 32250 24600 32310
rect 29760 32250 30120 32310
rect 33870 32250 34440 32310
rect 35310 32250 35880 32310
rect 36750 32250 37410 32310
rect 38280 32250 38760 32310
rect 39630 32250 39960 32310
rect 41160 32250 41400 32310
rect 42270 32250 42840 32310
rect 47160 32250 47490 32310
rect 49800 32250 50310 32310
rect 5130 26250 5520 26310
rect 14760 26250 15120 26310
rect 16110 26250 16530 26310
rect 17400 26250 17880 26310
rect 18750 26250 19080 26310
rect 20280 26250 20760 26310
rect 21630 26250 21960 26310
rect 22830 26250 23280 26310
rect 24270 26250 24840 26310
rect 27150 26250 28080 26310
rect 29400 26250 30210 26310
rect 35550 26250 35880 26310
rect 36750 26250 37410 26310
rect 38280 26250 38520 26310
rect 42270 26250 42840 26310
rect 44040 26250 44280 26310
rect 45480 26250 45720 26310
rect 50280 26250 50310 26310
rect 5130 20250 5160 20310
rect 7080 20250 8040 20310
rect 8910 20250 9120 20310
rect 10350 20250 10920 20310
rect 16080 20250 16680 20310
rect 17400 20250 17880 20310
rect 23160 20250 23760 20310
rect 27360 20250 27720 20310
rect 29790 20250 30120 20310
rect 31320 20250 31800 20310
rect 32670 20250 33000 20310
rect 33870 20250 34440 20310
rect 35310 20250 35640 20310
rect 39960 20250 40200 20310
rect 41070 20250 41400 20310
rect 42600 20250 43020 20310
rect 48120 20250 48600 20310
rect 49980 20250 50310 20310
rect 5130 14250 6120 14310
rect 6990 14250 7050 14310
rect 7200 14250 7560 14310
rect 12840 14250 13080 14310
rect 21720 14250 21960 14310
rect 23280 14250 23400 14310
rect 24270 14250 24690 14310
rect 27480 14250 27720 14310
rect 28590 14250 28920 14310
rect 35310 14250 35880 14310
rect 37080 14250 37560 14310
rect 40800 14250 41400 14310
rect 43320 14250 43440 14310
rect 43590 14250 44280 14310
rect 45480 14250 45960 14310
rect 46830 14250 47490 14310
rect 48360 14250 48840 14310
rect 50040 14250 50310 14310
rect 5130 8250 5400 8310
rect 12120 8250 12480 8310
rect 12630 8250 13560 8310
rect 15480 8250 15600 8310
rect 15840 8250 16200 8310
rect 24510 8250 25320 8310
rect 27240 8250 27720 8310
rect 28590 8250 29160 8310
rect 35040 8250 35490 8310
rect 39960 8250 40200 8310
rect 41070 8250 41400 8310
rect 44280 8250 44700 8310
rect 46920 8250 47490 8310
rect 48360 8250 48930 8310
rect 49800 8250 50310 8310
<< nwell >>
rect 5040 39540 50400 42660
rect 5040 33540 50400 36660
rect 5040 28950 50400 30660
rect 5040 27540 50220 28950
rect 5040 21540 50400 24660
rect 5040 15540 50400 18660
rect 5040 9540 50400 12660
rect 5040 4950 50400 6660
<< pwell >>
rect 5130 44100 44790 44250
rect 45450 44100 50310 44250
rect 5130 43950 50310 44100
rect 5400 43440 11640 43950
rect 12120 43440 13080 43950
rect 5400 43140 10680 43440
rect 13560 43140 14760 43950
rect 15240 43140 16110 43950
rect 16920 43140 18120 43950
rect 19080 43440 21720 43950
rect 19080 43140 21000 43440
rect 22440 43140 24360 43950
rect 24840 43140 26040 43950
rect 26520 43140 27390 43950
rect 27720 43140 29790 43950
rect 30120 43140 31320 43950
rect 31560 43140 32760 43950
rect 33090 43140 33960 43950
rect 34440 43440 35400 43950
rect 35640 43140 38760 43950
rect 39240 43140 41160 43950
rect 41640 43440 42360 43950
rect 42840 43440 49080 43950
rect 42840 43140 45240 43440
rect 45480 43140 49080 43440
rect 5730 38760 6600 39060
rect 5730 38250 6840 38760
rect 8130 38250 9000 39060
rect 9480 38760 10350 39060
rect 10680 38760 14190 39060
rect 14610 38760 15480 39060
rect 16200 38760 18600 39060
rect 19080 38760 20280 39060
rect 9480 38250 20280 38760
rect 20850 38760 23640 39060
rect 24600 38760 25800 39060
rect 20850 38250 25800 38760
rect 26100 38250 27480 39060
rect 27720 38250 28440 38760
rect 30450 38250 31320 39060
rect 31890 38250 32760 39060
rect 33240 38250 35160 39060
rect 35880 38250 37080 39060
rect 37650 38250 38520 39060
rect 38760 38250 39960 39060
rect 40200 38250 41070 39060
rect 41640 38250 42360 38760
rect 42840 38250 44040 39060
rect 44520 38250 45240 38760
rect 45720 38250 46920 39060
rect 47400 38250 48600 39060
rect 49170 38250 50040 39060
rect 5130 37950 50310 38250
rect 5490 37140 6360 37950
rect 6840 37440 7560 37950
rect 8040 37140 9240 37950
rect 10680 37140 11550 37950
rect 11880 37140 13080 37950
rect 14760 37140 15960 37950
rect 16530 37440 17640 37950
rect 16770 37140 17640 37440
rect 17880 37140 18750 37950
rect 19320 37140 20190 37950
rect 20760 37140 21630 37950
rect 22200 37140 23070 37950
rect 23640 37440 24360 37950
rect 24930 37140 25800 37950
rect 26280 37140 27480 37950
rect 27720 37140 28590 37950
rect 28920 37440 33960 37950
rect 28920 37140 31080 37440
rect 31800 37140 33960 37440
rect 34440 37140 37320 37950
rect 38760 37440 39480 37950
rect 39720 37140 41100 37950
rect 41400 37440 44040 37950
rect 42120 37140 43320 37440
rect 44280 37140 45480 37950
rect 45960 37140 46830 37950
rect 47400 37140 48600 37950
rect 49170 37140 50040 37950
rect 6360 32250 10680 33060
rect 10920 32250 12840 33060
rect 13560 32250 14280 32760
rect 15000 32250 15870 33060
rect 16440 32250 17640 33060
rect 19170 32250 20040 33060
rect 20850 32760 21720 33060
rect 20610 32250 21720 32760
rect 23160 32250 24360 33060
rect 24600 32250 27720 33060
rect 30930 32760 33870 33060
rect 30120 32250 33870 32760
rect 34440 32250 35310 33060
rect 35880 32250 36750 33060
rect 37410 32250 38280 33060
rect 38760 32250 39630 33060
rect 39960 32250 41160 33060
rect 41400 32250 42270 33060
rect 42840 32250 47160 33060
rect 47490 32250 48360 33060
rect 48930 32250 49800 33060
rect 5130 31950 50310 32250
rect 5160 31140 7080 31950
rect 7800 31140 9000 31950
rect 9570 31140 10440 31950
rect 10920 31140 12840 31950
rect 14520 31140 16440 31950
rect 16920 31140 18840 31950
rect 19080 31140 23160 31950
rect 23640 31440 24360 31950
rect 24690 31440 30120 31950
rect 24930 31140 27000 31440
rect 27570 31140 28440 31440
rect 28920 31140 30120 31440
rect 30600 31140 32520 31950
rect 33000 31140 33870 31950
rect 34440 31140 35310 31950
rect 35880 31140 37080 31950
rect 37560 31140 38430 31950
rect 38760 31140 39960 31950
rect 40440 31440 41160 31950
rect 41490 31140 42360 31950
rect 42840 31140 44040 31950
rect 44280 31140 45480 31950
rect 46050 31140 46920 31950
rect 47880 31140 49800 31950
rect 6840 26760 13470 27060
rect 13890 26760 14760 27060
rect 6840 26250 14760 26760
rect 15240 26250 16110 27060
rect 16530 26250 17400 27060
rect 17880 26250 18750 27060
rect 19080 26250 20280 27060
rect 20760 26250 21630 27060
rect 21960 26250 22830 27060
rect 23400 26250 24270 27060
rect 24840 26250 25710 27060
rect 26280 26250 27150 27060
rect 28200 26250 29400 27060
rect 30210 26250 31080 27060
rect 31560 26250 35550 27060
rect 35880 26250 36750 27060
rect 37410 26250 38280 27060
rect 38520 26250 42270 27060
rect 42840 26250 44040 27060
rect 44280 26250 45480 27060
rect 45720 26760 46920 27060
rect 47160 26760 50280 27060
rect 45720 26250 50280 26760
rect 5130 25950 50310 26250
rect 5160 25140 11160 25950
rect 11880 25440 12990 25950
rect 13560 25440 14280 25950
rect 12120 25140 12990 25440
rect 14760 25140 15960 25950
rect 20610 25140 21480 25950
rect 22920 25140 23790 25950
rect 25320 25140 27240 25950
rect 27720 25140 28920 25950
rect 30120 25440 32760 25950
rect 30840 25140 32040 25440
rect 33000 25140 33870 25950
rect 34440 25140 35310 25950
rect 35880 25140 36750 25950
rect 37320 25140 38190 25950
rect 38760 25140 39630 25950
rect 40200 25140 41070 25950
rect 41640 25140 42510 25950
rect 43080 25440 44040 25950
rect 44280 25440 45000 25950
rect 44520 25410 45000 25440
rect 47640 25140 49560 25950
rect 5160 20250 7080 21060
rect 8040 20250 8910 21060
rect 9480 20250 10350 21060
rect 10920 20250 12120 21060
rect 14040 20250 15960 21060
rect 16680 20250 17400 20760
rect 17880 20250 23160 21060
rect 24840 20250 25560 20760
rect 26040 20250 27240 21060
rect 27720 20250 29790 21060
rect 30120 20250 31320 21060
rect 31800 20250 32670 21060
rect 33000 20250 33870 21060
rect 34440 20250 35310 21060
rect 35640 20250 38520 21060
rect 38760 20250 39960 21060
rect 40200 20250 41070 21060
rect 41400 20250 42600 21060
rect 44040 20760 47640 21060
rect 43080 20250 48120 20760
rect 48600 20250 49980 21060
rect 5130 19950 50310 20250
rect 5400 19140 6600 19950
rect 8760 19140 10680 19950
rect 11400 19440 16440 19950
rect 11400 19140 16200 19440
rect 17640 19140 18840 19950
rect 19320 19140 20190 19950
rect 20760 19140 21630 19950
rect 21960 19140 22830 19950
rect 23400 19440 27720 19950
rect 23400 19140 27240 19440
rect 28200 19140 29400 19950
rect 30360 19140 31230 19950
rect 31800 19140 32670 19950
rect 33000 19140 34200 19950
rect 35640 19440 39630 19950
rect 35640 19140 36510 19440
rect 36840 19140 39630 19440
rect 40200 19140 41070 19950
rect 41400 19440 42120 19950
rect 42660 19140 44040 19950
rect 44280 19140 45480 19950
rect 45960 19140 46830 19950
rect 47400 19440 48360 19950
rect 48840 19140 50040 19950
rect 6120 14250 6990 15060
rect 7560 14250 12840 15060
rect 13080 14760 17400 15060
rect 17880 14760 19950 15060
rect 13080 14250 19950 14760
rect 20520 14250 21720 15060
rect 21960 14250 23160 15060
rect 23400 14250 24270 15060
rect 24690 14250 27480 15060
rect 27720 14250 28590 15060
rect 28920 14250 29790 15060
rect 30120 14250 33870 15060
rect 34440 14250 35310 15060
rect 35880 14250 37080 15060
rect 37560 14250 40440 15060
rect 41400 14250 43320 15060
rect 44280 14250 45480 15060
rect 45960 14250 46830 15060
rect 47490 14250 48360 15060
rect 48840 14250 50040 15060
rect 5130 13950 50310 14250
rect 6690 13140 7560 13950
rect 8760 13140 10200 13950
rect 10680 13140 11550 13950
rect 11880 13140 13080 13950
rect 15720 13140 21000 13950
rect 21720 13140 23640 13950
rect 24840 13140 26040 13950
rect 26520 13140 27390 13950
rect 28920 13140 31320 13950
rect 31890 13140 35640 13950
rect 35880 13140 36750 13950
rect 37320 13140 38190 13950
rect 38760 13140 39630 13950
rect 39960 13140 41160 13950
rect 41400 13440 42510 13950
rect 41400 13140 42270 13440
rect 43080 13140 43950 13950
rect 44280 13140 45480 13950
rect 45960 13140 46830 13950
rect 47400 13140 48600 13950
rect 49170 13140 50040 13950
rect 5400 8760 9480 9060
rect 9810 8760 10680 9060
rect 5400 8250 10680 8760
rect 11250 8250 12120 9060
rect 13560 8250 15480 9060
rect 16200 8250 24510 9060
rect 25320 8250 27240 9060
rect 27720 8250 28590 9060
rect 29160 8250 29880 8760
rect 30360 8250 31080 8760
rect 31560 8250 32760 9060
rect 33000 8250 34920 9060
rect 35730 8760 37470 9060
rect 37890 8760 39960 9060
rect 35490 8250 39960 8760
rect 40200 8250 41070 9060
rect 41400 8250 44280 9060
rect 45000 8250 46920 9060
rect 47490 8250 48360 9060
rect 48930 8250 49800 9060
rect 5130 7950 50310 8250
rect 5400 7140 7320 7950
rect 7800 7440 11880 7950
rect 8520 7140 11880 7440
rect 12120 7140 12990 7950
rect 13650 7440 14760 7950
rect 15240 7440 16200 7950
rect 17880 7440 18840 7950
rect 13650 7140 14520 7440
rect 20520 7140 21390 7950
rect 23160 7140 24030 7950
rect 25560 7140 27480 7950
rect 27720 7140 28590 7950
rect 28920 7140 33870 7950
rect 34530 7140 35400 7950
rect 35880 7140 36750 7950
rect 37320 7140 38520 7950
rect 38760 7140 39630 7950
rect 40200 7140 41070 7950
rect 43080 7440 44040 7950
rect 44340 7140 45720 7950
rect 46200 7440 46920 7950
rect 47160 7140 48360 7950
<< ntransistor >>
rect 5730 43320 5790 43920
rect 5970 43320 6030 43920
rect 6210 43320 6270 43920
rect 6930 43320 6990 43920
rect 7080 43320 7140 43920
rect 7890 43320 7950 43920
rect 8130 43320 8190 43920
rect 8370 43320 8430 43920
rect 9090 43320 9150 43920
rect 9360 43320 9420 43920
rect 9510 43320 9570 43920
rect 9870 43320 9930 43920
rect 10020 43320 10080 43920
rect 10290 43320 10350 43920
rect 11010 43620 11070 43920
rect 11250 43620 11310 43920
rect 12450 43620 12510 43920
rect 12690 43620 12750 43920
rect 13890 43320 13950 43920
rect 14130 43320 14190 43920
rect 14370 43320 14430 43920
rect 15570 43320 15630 43920
rect 15720 43320 15780 43920
rect 17250 43320 17310 43920
rect 17490 43320 17550 43920
rect 17730 43320 17790 43920
rect 19410 43320 19470 43920
rect 19680 43320 19740 43920
rect 19830 43320 19890 43920
rect 20190 43320 20250 43920
rect 20340 43320 20400 43920
rect 20610 43320 20670 43920
rect 21330 43620 21390 43920
rect 22770 43320 22830 43920
rect 23040 43320 23100 43920
rect 23190 43320 23250 43920
rect 23550 43320 23610 43920
rect 23700 43320 23760 43920
rect 23970 43320 24030 43920
rect 25170 43320 25230 43920
rect 25410 43320 25470 43920
rect 25650 43320 25710 43920
rect 26850 43320 26910 43920
rect 27000 43320 27060 43920
rect 28050 43320 28110 43920
rect 28290 43320 28350 43920
rect 28530 43320 28590 43920
rect 29250 43320 29310 43920
rect 29400 43320 29460 43920
rect 30450 43320 30510 43920
rect 30690 43320 30750 43920
rect 30930 43320 30990 43920
rect 31890 43320 31950 43920
rect 32130 43320 32190 43920
rect 32370 43320 32430 43920
rect 33420 43320 33480 43920
rect 33570 43320 33630 43920
rect 34770 43620 34830 43920
rect 35010 43620 35070 43920
rect 35970 43320 36030 43920
rect 36240 43320 36300 43920
rect 36390 43320 36450 43920
rect 36750 43320 36810 43920
rect 36900 43320 36960 43920
rect 37170 43320 37230 43920
rect 37890 43320 37950 43920
rect 38130 43320 38190 43920
rect 38370 43320 38430 43920
rect 39570 43320 39630 43920
rect 39840 43320 39900 43920
rect 39990 43320 40050 43920
rect 40350 43320 40410 43920
rect 40500 43320 40560 43920
rect 40770 43320 40830 43920
rect 41970 43620 42030 43920
rect 43170 43320 43230 43920
rect 43410 43320 43470 43920
rect 43650 43320 43710 43920
rect 44370 43320 44430 43920
rect 44610 43320 44670 43920
rect 44850 43320 44910 43920
rect 45330 43620 45390 43920
rect 45810 43320 45870 43920
rect 46080 43320 46140 43920
rect 46230 43320 46290 43920
rect 46590 43320 46650 43920
rect 46740 43320 46800 43920
rect 47010 43320 47070 43920
rect 47490 43320 47550 43920
rect 47760 43320 47820 43920
rect 47910 43320 47970 43920
rect 48270 43320 48330 43920
rect 48420 43320 48480 43920
rect 48690 43320 48750 43920
rect 6060 38280 6120 38880
rect 6210 38280 6270 38880
rect 6450 38280 6510 38580
rect 8460 38280 8520 38880
rect 8610 38280 8670 38880
rect 9810 38280 9870 38880
rect 9960 38280 10020 38880
rect 10770 38280 10830 38580
rect 11010 38280 11070 38880
rect 11160 38280 11220 38880
rect 11730 38280 11790 38880
rect 12000 38280 12060 38880
rect 12150 38280 12210 38880
rect 12510 38280 12570 38880
rect 12660 38280 12720 38880
rect 12930 38280 12990 38880
rect 13650 38280 13710 38880
rect 13800 38280 13860 38880
rect 14700 38280 14760 38580
rect 14940 38280 15000 38880
rect 15090 38280 15150 38880
rect 15810 38280 15870 38580
rect 16530 38280 16590 38880
rect 16770 38280 16830 38880
rect 17010 38280 17070 38880
rect 17730 38280 17790 38880
rect 17970 38280 18030 38880
rect 18210 38280 18270 38880
rect 18690 38280 18750 38580
rect 19410 38280 19470 38880
rect 19650 38280 19710 38880
rect 19890 38280 19950 38880
rect 21180 38280 21240 38880
rect 21330 38280 21390 38880
rect 22050 38280 22110 38880
rect 22320 38280 22380 38880
rect 22470 38280 22530 38880
rect 22830 38280 22890 38880
rect 22980 38280 23040 38880
rect 23250 38280 23310 38880
rect 23970 38280 24030 38580
rect 24210 38280 24270 38580
rect 24930 38280 24990 38880
rect 25170 38280 25230 38880
rect 25410 38280 25470 38880
rect 26430 38280 26490 38880
rect 26580 38280 26640 38880
rect 26940 38280 27000 38880
rect 27090 38280 27150 38880
rect 28050 38280 28110 38580
rect 30780 38280 30840 38880
rect 30930 38280 30990 38880
rect 32220 38280 32280 38880
rect 32370 38280 32430 38880
rect 33570 38280 33630 38880
rect 33840 38280 33900 38880
rect 33990 38280 34050 38880
rect 34350 38280 34410 38880
rect 34500 38280 34560 38880
rect 34770 38280 34830 38880
rect 36210 38280 36270 38880
rect 36450 38280 36510 38880
rect 36690 38280 36750 38880
rect 37980 38280 38040 38880
rect 38130 38280 38190 38880
rect 39090 38280 39150 38880
rect 39330 38280 39390 38880
rect 39570 38280 39630 38880
rect 40530 38280 40590 38880
rect 40680 38280 40740 38880
rect 41970 38280 42030 38580
rect 43170 38280 43230 38880
rect 43410 38280 43470 38880
rect 43650 38280 43710 38880
rect 44850 38280 44910 38580
rect 46050 38280 46110 38880
rect 46290 38280 46350 38880
rect 46530 38280 46590 38880
rect 47730 38280 47790 38880
rect 47970 38280 48030 38880
rect 48210 38280 48270 38880
rect 49500 38280 49560 38880
rect 49650 38280 49710 38880
rect 5820 37320 5880 37920
rect 5970 37320 6030 37920
rect 7170 37620 7230 37920
rect 8370 37320 8430 37920
rect 8610 37320 8670 37920
rect 8850 37320 8910 37920
rect 11010 37320 11070 37920
rect 11160 37320 11220 37920
rect 12210 37320 12270 37920
rect 12450 37320 12510 37920
rect 12690 37320 12750 37920
rect 15090 37320 15150 37920
rect 15330 37320 15390 37920
rect 15570 37320 15630 37920
rect 16860 37620 16920 37920
rect 17100 37320 17160 37920
rect 17250 37320 17310 37920
rect 18210 37320 18270 37920
rect 18360 37320 18420 37920
rect 19650 37320 19710 37920
rect 19800 37320 19860 37920
rect 21090 37320 21150 37920
rect 21240 37320 21300 37920
rect 22530 37320 22590 37920
rect 22680 37320 22740 37920
rect 23970 37620 24030 37920
rect 25260 37320 25320 37920
rect 25410 37320 25470 37920
rect 26610 37320 26670 37920
rect 26850 37320 26910 37920
rect 27090 37320 27150 37920
rect 28050 37320 28110 37920
rect 28200 37320 28260 37920
rect 29250 37320 29310 37920
rect 29400 37320 29460 37920
rect 30210 37320 30270 37920
rect 30450 37320 30510 37920
rect 30690 37320 30750 37920
rect 31410 37620 31470 37920
rect 32130 37320 32190 37920
rect 32370 37320 32430 37920
rect 32610 37320 32670 37920
rect 33420 37320 33480 37920
rect 33570 37320 33630 37920
rect 34770 37320 34830 37920
rect 34920 37320 34980 37920
rect 35730 37320 35790 37920
rect 36000 37320 36060 37920
rect 36150 37320 36210 37920
rect 36510 37320 36570 37920
rect 36660 37320 36720 37920
rect 36930 37320 36990 37920
rect 39090 37620 39150 37920
rect 40050 37320 40110 37920
rect 40200 37320 40260 37920
rect 40560 37320 40620 37920
rect 40710 37320 40770 37920
rect 41730 37620 41790 37920
rect 42450 37320 42510 37920
rect 42690 37320 42750 37920
rect 42930 37320 42990 37920
rect 43650 37620 43710 37920
rect 44610 37320 44670 37920
rect 44850 37320 44910 37920
rect 45090 37320 45150 37920
rect 46290 37320 46350 37920
rect 46440 37320 46500 37920
rect 47730 37320 47790 37920
rect 47970 37320 48030 37920
rect 48210 37320 48270 37920
rect 49500 37320 49560 37920
rect 49650 37320 49710 37920
rect 6690 32280 6750 32880
rect 6930 32280 6990 32880
rect 7170 32280 7230 32880
rect 7890 32280 7950 32880
rect 8130 32280 8190 32880
rect 8370 32280 8430 32880
rect 9090 32280 9150 32880
rect 9360 32280 9420 32880
rect 9510 32280 9570 32880
rect 9870 32280 9930 32880
rect 10020 32280 10080 32880
rect 10290 32280 10350 32880
rect 11250 32280 11310 32880
rect 11520 32280 11580 32880
rect 11670 32280 11730 32880
rect 12030 32280 12090 32880
rect 12180 32280 12240 32880
rect 12450 32280 12510 32880
rect 13890 32280 13950 32580
rect 15330 32280 15390 32880
rect 15480 32280 15540 32880
rect 16770 32280 16830 32880
rect 17010 32280 17070 32880
rect 17250 32280 17310 32880
rect 19500 32280 19560 32880
rect 19650 32280 19710 32880
rect 20940 32280 21000 32580
rect 21180 32280 21240 32880
rect 21330 32280 21390 32880
rect 23490 32280 23550 32880
rect 23730 32280 23790 32880
rect 23970 32280 24030 32880
rect 24930 32280 24990 32880
rect 25170 32280 25230 32880
rect 25410 32280 25470 32880
rect 26130 32280 26190 32880
rect 26400 32280 26460 32880
rect 26550 32280 26610 32880
rect 26910 32280 26970 32880
rect 27060 32280 27120 32880
rect 27330 32280 27390 32880
rect 30450 32280 30510 32580
rect 31260 32280 31320 32880
rect 31410 32280 31470 32880
rect 32130 32280 32190 32880
rect 32370 32280 32430 32880
rect 32610 32280 32670 32880
rect 33330 32280 33390 32880
rect 33480 32280 33540 32880
rect 34770 32280 34830 32880
rect 34920 32280 34980 32880
rect 36210 32280 36270 32880
rect 36360 32280 36420 32880
rect 37740 32280 37800 32880
rect 37890 32280 37950 32880
rect 39090 32280 39150 32880
rect 39240 32280 39300 32880
rect 40290 32280 40350 32880
rect 40530 32280 40590 32880
rect 40770 32280 40830 32880
rect 41730 32280 41790 32880
rect 41880 32280 41940 32880
rect 43170 32280 43230 32880
rect 43410 32280 43470 32880
rect 43650 32280 43710 32880
rect 44370 32280 44430 32880
rect 44640 32280 44700 32880
rect 44790 32280 44850 32880
rect 45150 32280 45210 32880
rect 45300 32280 45360 32880
rect 45570 32280 45630 32880
rect 46290 32280 46350 32880
rect 46530 32280 46590 32880
rect 46770 32280 46830 32880
rect 47820 32280 47880 32880
rect 47970 32280 48030 32880
rect 49260 32280 49320 32880
rect 49410 32280 49470 32880
rect 5490 31320 5550 31920
rect 5760 31320 5820 31920
rect 5910 31320 5970 31920
rect 6270 31320 6330 31920
rect 6420 31320 6480 31920
rect 6690 31320 6750 31920
rect 8130 31320 8190 31920
rect 8370 31320 8430 31920
rect 8610 31320 8670 31920
rect 9900 31320 9960 31920
rect 10050 31320 10110 31920
rect 11250 31320 11310 31920
rect 11520 31320 11580 31920
rect 11670 31320 11730 31920
rect 12030 31320 12090 31920
rect 12180 31320 12240 31920
rect 12450 31320 12510 31920
rect 14850 31320 14910 31920
rect 15120 31320 15180 31920
rect 15270 31320 15330 31920
rect 15630 31320 15690 31920
rect 15780 31320 15840 31920
rect 16050 31320 16110 31920
rect 17250 31320 17310 31920
rect 17520 31320 17580 31920
rect 17670 31320 17730 31920
rect 18030 31320 18090 31920
rect 18180 31320 18240 31920
rect 18450 31320 18510 31920
rect 19410 31320 19470 31920
rect 19680 31320 19740 31920
rect 19830 31320 19890 31920
rect 20190 31320 20250 31920
rect 20340 31320 20400 31920
rect 20610 31320 20670 31920
rect 21330 31320 21390 31920
rect 21480 31320 21540 31920
rect 22290 31320 22350 31920
rect 22530 31320 22590 31920
rect 22770 31320 22830 31920
rect 23970 31620 24030 31920
rect 25020 31620 25080 31920
rect 25260 31320 25320 31920
rect 25410 31320 25470 31920
rect 26130 31320 26190 31920
rect 26370 31320 26430 31920
rect 26610 31320 26670 31920
rect 27330 31620 27390 31920
rect 27900 31320 27960 31920
rect 28050 31320 28110 31920
rect 28770 31620 28830 31920
rect 29250 31320 29310 31920
rect 29490 31320 29550 31920
rect 29730 31320 29790 31920
rect 30930 31320 30990 31920
rect 31200 31320 31260 31920
rect 31350 31320 31410 31920
rect 31710 31320 31770 31920
rect 31860 31320 31920 31920
rect 32130 31320 32190 31920
rect 33330 31320 33390 31920
rect 33480 31320 33540 31920
rect 34770 31320 34830 31920
rect 34920 31320 34980 31920
rect 36210 31320 36270 31920
rect 36450 31320 36510 31920
rect 36690 31320 36750 31920
rect 37890 31320 37950 31920
rect 38040 31320 38100 31920
rect 39090 31320 39150 31920
rect 39330 31320 39390 31920
rect 39570 31320 39630 31920
rect 40770 31620 40830 31920
rect 41820 31320 41880 31920
rect 41970 31320 42030 31920
rect 43170 31320 43230 31920
rect 43410 31320 43470 31920
rect 43650 31320 43710 31920
rect 44610 31320 44670 31920
rect 44850 31320 44910 31920
rect 45090 31320 45150 31920
rect 46380 31320 46440 31920
rect 46530 31320 46590 31920
rect 48210 31320 48270 31920
rect 48480 31320 48540 31920
rect 48630 31320 48690 31920
rect 48990 31320 49050 31920
rect 49140 31320 49200 31920
rect 49410 31320 49470 31920
rect 7170 26280 7230 26880
rect 7440 26280 7500 26880
rect 7590 26280 7650 26880
rect 7950 26280 8010 26880
rect 8100 26280 8160 26880
rect 8370 26280 8430 26880
rect 8850 26280 8910 26880
rect 9000 26280 9060 26880
rect 9570 26280 9630 26880
rect 9840 26280 9900 26880
rect 9990 26280 10050 26880
rect 10350 26280 10410 26880
rect 10500 26280 10560 26880
rect 10770 26280 10830 26880
rect 11250 26280 11310 26880
rect 11490 26280 11550 26880
rect 11730 26280 11790 26880
rect 12210 26280 12270 26880
rect 12360 26280 12420 26880
rect 12930 26280 12990 26880
rect 13080 26280 13140 26880
rect 13980 26280 14040 26580
rect 14220 26280 14280 26880
rect 14370 26280 14430 26880
rect 15570 26280 15630 26880
rect 15720 26280 15780 26880
rect 16860 26280 16920 26880
rect 17010 26280 17070 26880
rect 18210 26280 18270 26880
rect 18360 26280 18420 26880
rect 19410 26280 19470 26880
rect 19650 26280 19710 26880
rect 19890 26280 19950 26880
rect 21090 26280 21150 26880
rect 21240 26280 21300 26880
rect 22290 26280 22350 26880
rect 22440 26280 22500 26880
rect 23730 26280 23790 26880
rect 23880 26280 23940 26880
rect 25170 26280 25230 26880
rect 25320 26280 25380 26880
rect 26610 26280 26670 26880
rect 26760 26280 26820 26880
rect 28530 26280 28590 26880
rect 28770 26280 28830 26880
rect 29010 26280 29070 26880
rect 30540 26280 30600 26880
rect 30690 26280 30750 26880
rect 31890 26280 31950 26880
rect 32130 26280 32190 26880
rect 32370 26280 32430 26880
rect 33090 26280 33150 26880
rect 33360 26280 33420 26880
rect 33510 26280 33570 26880
rect 33870 26280 33930 26880
rect 34020 26280 34080 26880
rect 34290 26280 34350 26880
rect 35010 26280 35070 26880
rect 35160 26280 35220 26880
rect 36210 26280 36270 26880
rect 36360 26280 36420 26880
rect 37740 26280 37800 26880
rect 37890 26280 37950 26880
rect 38850 26280 38910 26880
rect 39000 26280 39060 26880
rect 39810 26280 39870 26880
rect 40080 26280 40140 26880
rect 40230 26280 40290 26880
rect 40590 26280 40650 26880
rect 40740 26280 40800 26880
rect 41010 26280 41070 26880
rect 41730 26280 41790 26880
rect 41880 26280 41940 26880
rect 43170 26280 43230 26880
rect 43410 26280 43470 26880
rect 43650 26280 43710 26880
rect 44610 26280 44670 26880
rect 44850 26280 44910 26880
rect 45090 26280 45150 26880
rect 46050 26280 46110 26880
rect 46290 26280 46350 26880
rect 46530 26280 46590 26880
rect 47010 26280 47070 26580
rect 47490 26280 47550 26880
rect 47640 26280 47700 26880
rect 48000 26280 48060 26880
rect 48150 26280 48210 26880
rect 48690 26280 48750 26880
rect 48840 26280 48900 26880
rect 49410 26280 49470 26880
rect 49650 26280 49710 26880
rect 49890 26280 49950 26880
rect 5490 25320 5550 25920
rect 5760 25320 5820 25920
rect 5910 25320 5970 25920
rect 6270 25320 6330 25920
rect 6420 25320 6480 25920
rect 6690 25320 6750 25920
rect 7170 25320 7230 25920
rect 7320 25320 7380 25920
rect 7890 25320 7950 25920
rect 8130 25320 8190 25920
rect 8370 25320 8430 25920
rect 8850 25320 8910 25920
rect 9000 25320 9060 25920
rect 9570 25320 9630 25920
rect 9840 25320 9900 25920
rect 9990 25320 10050 25920
rect 10350 25320 10410 25920
rect 10500 25320 10560 25920
rect 10770 25320 10830 25920
rect 12210 25620 12270 25920
rect 12450 25320 12510 25920
rect 12600 25320 12660 25920
rect 13890 25620 13950 25920
rect 15090 25320 15150 25920
rect 15330 25320 15390 25920
rect 15570 25320 15630 25920
rect 20940 25320 21000 25920
rect 21090 25320 21150 25920
rect 23250 25320 23310 25920
rect 23400 25320 23460 25920
rect 25650 25320 25710 25920
rect 25920 25320 25980 25920
rect 26070 25320 26130 25920
rect 26430 25320 26490 25920
rect 26580 25320 26640 25920
rect 26850 25320 26910 25920
rect 28050 25320 28110 25920
rect 28290 25320 28350 25920
rect 28530 25320 28590 25920
rect 30450 25620 30510 25920
rect 31170 25320 31230 25920
rect 31410 25320 31470 25920
rect 31650 25320 31710 25920
rect 32370 25620 32430 25920
rect 33330 25320 33390 25920
rect 33480 25320 33540 25920
rect 34770 25320 34830 25920
rect 34920 25320 34980 25920
rect 36210 25320 36270 25920
rect 36360 25320 36420 25920
rect 37650 25320 37710 25920
rect 37800 25320 37860 25920
rect 39090 25320 39150 25920
rect 39240 25320 39300 25920
rect 40530 25320 40590 25920
rect 40680 25320 40740 25920
rect 41970 25320 42030 25920
rect 42120 25320 42180 25920
rect 43410 25620 43470 25920
rect 43650 25620 43710 25920
rect 44610 25620 44670 25920
rect 47970 25320 48030 25920
rect 48240 25320 48300 25920
rect 48390 25320 48450 25920
rect 48750 25320 48810 25920
rect 48900 25320 48960 25920
rect 49170 25320 49230 25920
rect 5490 20280 5550 20880
rect 5760 20280 5820 20880
rect 5910 20280 5970 20880
rect 6270 20280 6330 20880
rect 6420 20280 6480 20880
rect 6690 20280 6750 20880
rect 8370 20280 8430 20880
rect 8520 20280 8580 20880
rect 9810 20280 9870 20880
rect 9960 20280 10020 20880
rect 11250 20280 11310 20880
rect 11490 20280 11550 20880
rect 11730 20280 11790 20880
rect 14370 20280 14430 20880
rect 14640 20280 14700 20880
rect 14790 20280 14850 20880
rect 15150 20280 15210 20880
rect 15300 20280 15360 20880
rect 15570 20280 15630 20880
rect 17010 20280 17070 20580
rect 18210 20280 18270 20880
rect 18360 20280 18420 20880
rect 18930 20280 18990 20880
rect 19200 20280 19260 20880
rect 19350 20280 19410 20880
rect 19710 20280 19770 20880
rect 19860 20280 19920 20880
rect 20130 20280 20190 20880
rect 20610 20280 20670 20880
rect 20880 20280 20940 20880
rect 21030 20280 21090 20880
rect 21390 20280 21450 20880
rect 21540 20280 21600 20880
rect 21810 20280 21870 20880
rect 22290 20280 22350 20880
rect 22530 20280 22590 20880
rect 22770 20280 22830 20880
rect 25170 20280 25230 20580
rect 26370 20280 26430 20880
rect 26610 20280 26670 20880
rect 26850 20280 26910 20880
rect 28050 20280 28110 20880
rect 28290 20280 28350 20880
rect 28530 20280 28590 20880
rect 29250 20280 29310 20880
rect 29400 20280 29460 20880
rect 30450 20280 30510 20880
rect 30690 20280 30750 20880
rect 30930 20280 30990 20880
rect 32130 20280 32190 20880
rect 32280 20280 32340 20880
rect 33330 20280 33390 20880
rect 33480 20280 33540 20880
rect 34770 20280 34830 20880
rect 34920 20280 34980 20880
rect 35970 20280 36030 20880
rect 36120 20280 36180 20880
rect 36930 20280 36990 20880
rect 37200 20280 37260 20880
rect 37350 20280 37410 20880
rect 37710 20280 37770 20880
rect 37860 20280 37920 20880
rect 38130 20280 38190 20880
rect 39090 20280 39150 20880
rect 39330 20280 39390 20880
rect 39570 20280 39630 20880
rect 40530 20280 40590 20880
rect 40680 20280 40740 20880
rect 41730 20280 41790 20880
rect 41970 20280 42030 20880
rect 42210 20280 42270 20880
rect 43410 20280 43470 20580
rect 43650 20280 43710 20580
rect 44370 20280 44430 20880
rect 44640 20280 44700 20880
rect 44790 20280 44850 20880
rect 45150 20280 45210 20880
rect 45300 20280 45360 20880
rect 45570 20280 45630 20880
rect 46050 20280 46110 20880
rect 46320 20280 46380 20880
rect 46470 20280 46530 20880
rect 46830 20280 46890 20880
rect 46980 20280 47040 20880
rect 47250 20280 47310 20880
rect 47730 20280 47790 20580
rect 48930 20280 48990 20880
rect 49080 20280 49140 20880
rect 49440 20280 49500 20880
rect 49590 20280 49650 20880
rect 5730 19320 5790 19920
rect 5970 19320 6030 19920
rect 6210 19320 6270 19920
rect 9090 19320 9150 19920
rect 9360 19320 9420 19920
rect 9510 19320 9570 19920
rect 9870 19320 9930 19920
rect 10020 19320 10080 19920
rect 10290 19320 10350 19920
rect 11730 19320 11790 19920
rect 12000 19320 12060 19920
rect 12150 19320 12210 19920
rect 12510 19320 12570 19920
rect 12660 19320 12720 19920
rect 12930 19320 12990 19920
rect 13650 19320 13710 19920
rect 13920 19320 13980 19920
rect 14070 19320 14130 19920
rect 14430 19320 14490 19920
rect 14580 19320 14640 19920
rect 14850 19320 14910 19920
rect 15660 19320 15720 19920
rect 15810 19320 15870 19920
rect 16050 19620 16110 19920
rect 17970 19320 18030 19920
rect 18210 19320 18270 19920
rect 18450 19320 18510 19920
rect 19650 19320 19710 19920
rect 19800 19320 19860 19920
rect 21090 19320 21150 19920
rect 21240 19320 21300 19920
rect 22290 19320 22350 19920
rect 22440 19320 22500 19920
rect 23730 19320 23790 19920
rect 23880 19320 23940 19920
rect 24690 19320 24750 19920
rect 24960 19320 25020 19920
rect 25110 19320 25170 19920
rect 25470 19320 25530 19920
rect 25620 19320 25680 19920
rect 25890 19320 25950 19920
rect 26370 19320 26430 19920
rect 26610 19320 26670 19920
rect 26850 19320 26910 19920
rect 27330 19620 27390 19920
rect 28530 19320 28590 19920
rect 28770 19320 28830 19920
rect 29010 19320 29070 19920
rect 30690 19320 30750 19920
rect 30840 19320 30900 19920
rect 32130 19320 32190 19920
rect 32280 19320 32340 19920
rect 33330 19320 33390 19920
rect 33570 19320 33630 19920
rect 33810 19320 33870 19920
rect 35970 19320 36030 19920
rect 36120 19320 36180 19920
rect 36930 19620 36990 19920
rect 37170 19320 37230 19920
rect 37320 19320 37380 19920
rect 38130 19320 38190 19920
rect 38280 19320 38340 19920
rect 39090 19320 39150 19920
rect 39240 19320 39300 19920
rect 40530 19320 40590 19920
rect 40680 19320 40740 19920
rect 41730 19620 41790 19920
rect 42990 19320 43050 19920
rect 43140 19320 43200 19920
rect 43500 19320 43560 19920
rect 43650 19320 43710 19920
rect 44610 19320 44670 19920
rect 44850 19320 44910 19920
rect 45090 19320 45150 19920
rect 46290 19320 46350 19920
rect 46440 19320 46500 19920
rect 47730 19620 47790 19920
rect 47970 19620 48030 19920
rect 49170 19320 49230 19920
rect 49410 19320 49470 19920
rect 49650 19320 49710 19920
rect 6450 14280 6510 14880
rect 6600 14280 6660 14880
rect 7890 14280 7950 14880
rect 8160 14280 8220 14880
rect 8310 14280 8370 14880
rect 8670 14280 8730 14880
rect 8820 14280 8880 14880
rect 9090 14280 9150 14880
rect 9570 14280 9630 14880
rect 9840 14280 9900 14880
rect 9990 14280 10050 14880
rect 10350 14280 10410 14880
rect 10500 14280 10560 14880
rect 10770 14280 10830 14880
rect 11250 14280 11310 14880
rect 11520 14280 11580 14880
rect 11670 14280 11730 14880
rect 12030 14280 12090 14880
rect 12180 14280 12240 14880
rect 12450 14280 12510 14880
rect 13410 14280 13470 14880
rect 13680 14280 13740 14880
rect 13830 14280 13890 14880
rect 14190 14280 14250 14880
rect 14340 14280 14400 14880
rect 14610 14280 14670 14880
rect 15090 14280 15150 14880
rect 15360 14280 15420 14880
rect 15510 14280 15570 14880
rect 15870 14280 15930 14880
rect 16020 14280 16080 14880
rect 16290 14280 16350 14880
rect 16860 14280 16920 14880
rect 17010 14280 17070 14880
rect 17250 14280 17310 14580
rect 17730 14280 17790 14580
rect 18210 14280 18270 14880
rect 18450 14280 18510 14880
rect 18690 14280 18750 14880
rect 19410 14280 19470 14880
rect 19560 14280 19620 14880
rect 20850 14280 20910 14880
rect 21090 14280 21150 14880
rect 21330 14280 21390 14880
rect 22290 14280 22350 14880
rect 22530 14280 22590 14880
rect 22770 14280 22830 14880
rect 23730 14280 23790 14880
rect 23880 14280 23940 14880
rect 25020 14280 25080 14880
rect 25170 14280 25230 14880
rect 25890 14280 25950 14880
rect 26160 14280 26220 14880
rect 26310 14280 26370 14880
rect 26670 14280 26730 14880
rect 26820 14280 26880 14880
rect 27090 14280 27150 14880
rect 28050 14280 28110 14880
rect 28200 14280 28260 14880
rect 29250 14280 29310 14880
rect 29400 14280 29460 14880
rect 30450 14280 30510 14880
rect 30720 14280 30780 14880
rect 30870 14280 30930 14880
rect 31230 14280 31290 14880
rect 31380 14280 31440 14880
rect 31650 14280 31710 14880
rect 32460 14280 32520 14880
rect 32610 14280 32670 14880
rect 33330 14280 33390 14880
rect 33480 14280 33540 14880
rect 34770 14280 34830 14880
rect 34920 14280 34980 14880
rect 36210 14280 36270 14880
rect 36450 14280 36510 14880
rect 36690 14280 36750 14880
rect 37890 14280 37950 14880
rect 38040 14280 38100 14880
rect 38850 14280 38910 14880
rect 39120 14280 39180 14880
rect 39270 14280 39330 14880
rect 39630 14280 39690 14880
rect 39780 14280 39840 14880
rect 40050 14280 40110 14880
rect 41730 14280 41790 14880
rect 42000 14280 42060 14880
rect 42150 14280 42210 14880
rect 42510 14280 42570 14880
rect 42660 14280 42720 14880
rect 42930 14280 42990 14880
rect 44610 14280 44670 14880
rect 44850 14280 44910 14880
rect 45090 14280 45150 14880
rect 46290 14280 46350 14880
rect 46440 14280 46500 14880
rect 47820 14280 47880 14880
rect 47970 14280 48030 14880
rect 49170 14280 49230 14880
rect 49410 14280 49470 14880
rect 49650 14280 49710 14880
rect 7020 13320 7080 13920
rect 7170 13320 7230 13920
rect 9090 13320 9150 13920
rect 9330 13320 9390 13920
rect 9570 13320 9630 13920
rect 9810 13320 9870 13920
rect 11010 13320 11070 13920
rect 11160 13320 11220 13920
rect 12210 13320 12270 13920
rect 12450 13320 12510 13920
rect 12690 13320 12750 13920
rect 16050 13320 16110 13920
rect 16200 13320 16260 13920
rect 16770 13320 16830 13920
rect 17010 13320 17070 13920
rect 17250 13320 17310 13920
rect 17730 13320 17790 13920
rect 18000 13320 18060 13920
rect 18150 13320 18210 13920
rect 18510 13320 18570 13920
rect 18660 13320 18720 13920
rect 18930 13320 18990 13920
rect 19410 13320 19470 13920
rect 19680 13320 19740 13920
rect 19830 13320 19890 13920
rect 20190 13320 20250 13920
rect 20340 13320 20400 13920
rect 20610 13320 20670 13920
rect 22050 13320 22110 13920
rect 22320 13320 22380 13920
rect 22470 13320 22530 13920
rect 22830 13320 22890 13920
rect 22980 13320 23040 13920
rect 23250 13320 23310 13920
rect 25170 13320 25230 13920
rect 25410 13320 25470 13920
rect 25650 13320 25710 13920
rect 26850 13320 26910 13920
rect 27000 13320 27060 13920
rect 29250 13320 29310 13920
rect 29490 13320 29550 13920
rect 29730 13320 29790 13920
rect 30450 13320 30510 13920
rect 30690 13320 30750 13920
rect 30930 13320 30990 13920
rect 32220 13320 32280 13920
rect 32370 13320 32430 13920
rect 33090 13320 33150 13920
rect 33360 13320 33420 13920
rect 33510 13320 33570 13920
rect 33870 13320 33930 13920
rect 34020 13320 34080 13920
rect 34290 13320 34350 13920
rect 34770 13320 34830 13920
rect 35010 13320 35070 13920
rect 35250 13320 35310 13920
rect 36210 13320 36270 13920
rect 36360 13320 36420 13920
rect 37650 13320 37710 13920
rect 37800 13320 37860 13920
rect 39090 13320 39150 13920
rect 39240 13320 39300 13920
rect 40290 13320 40350 13920
rect 40530 13320 40590 13920
rect 40770 13320 40830 13920
rect 41730 13320 41790 13920
rect 41880 13320 41940 13920
rect 42120 13620 42180 13920
rect 43410 13320 43470 13920
rect 43560 13320 43620 13920
rect 44610 13320 44670 13920
rect 44850 13320 44910 13920
rect 45090 13320 45150 13920
rect 46290 13320 46350 13920
rect 46440 13320 46500 13920
rect 47730 13320 47790 13920
rect 47970 13320 48030 13920
rect 48210 13320 48270 13920
rect 49500 13320 49560 13920
rect 49650 13320 49710 13920
rect 5730 8280 5790 8880
rect 5970 8280 6030 8880
rect 6210 8280 6270 8880
rect 6930 8280 6990 8880
rect 7080 8280 7140 8880
rect 7890 8280 7950 8880
rect 8160 8280 8220 8880
rect 8310 8280 8370 8880
rect 8670 8280 8730 8880
rect 8820 8280 8880 8880
rect 9090 8280 9150 8880
rect 9900 8280 9960 8580
rect 10140 8280 10200 8880
rect 10290 8280 10350 8880
rect 11580 8280 11640 8880
rect 11730 8280 11790 8880
rect 13890 8280 13950 8880
rect 14160 8280 14220 8880
rect 14310 8280 14370 8880
rect 14670 8280 14730 8880
rect 14820 8280 14880 8880
rect 15090 8280 15150 8880
rect 16530 8280 16590 8880
rect 16680 8280 16740 8880
rect 17490 8280 17550 8880
rect 17760 8280 17820 8880
rect 17910 8280 17970 8880
rect 18270 8280 18330 8880
rect 18420 8280 18480 8880
rect 18690 8280 18750 8880
rect 19410 8280 19470 8880
rect 19680 8280 19740 8880
rect 19830 8280 19890 8880
rect 20190 8280 20250 8880
rect 20340 8280 20400 8880
rect 20610 8280 20670 8880
rect 21420 8280 21480 8880
rect 21570 8280 21630 8880
rect 22050 8280 22110 8880
rect 22320 8280 22380 8880
rect 22470 8280 22530 8880
rect 22830 8280 22890 8880
rect 22980 8280 23040 8880
rect 23250 8280 23310 8880
rect 23970 8280 24030 8880
rect 24120 8280 24180 8880
rect 25650 8280 25710 8880
rect 25920 8280 25980 8880
rect 26070 8280 26130 8880
rect 26430 8280 26490 8880
rect 26580 8280 26640 8880
rect 26850 8280 26910 8880
rect 28050 8280 28110 8880
rect 28200 8280 28260 8880
rect 29490 8280 29550 8580
rect 30690 8280 30750 8580
rect 31890 8280 31950 8880
rect 32130 8280 32190 8880
rect 32370 8280 32430 8880
rect 33330 8280 33390 8880
rect 33600 8280 33660 8880
rect 33750 8280 33810 8880
rect 34110 8280 34170 8880
rect 34260 8280 34320 8880
rect 34530 8280 34590 8880
rect 35820 8280 35880 8580
rect 36060 8280 36120 8880
rect 36210 8280 36270 8880
rect 36930 8280 36990 8880
rect 37080 8280 37140 8880
rect 37980 8280 38040 8580
rect 38220 8280 38280 8880
rect 38370 8280 38430 8880
rect 39090 8280 39150 8880
rect 39330 8280 39390 8880
rect 39570 8280 39630 8880
rect 40530 8280 40590 8880
rect 40680 8280 40740 8880
rect 41730 8280 41790 8880
rect 41880 8280 41940 8880
rect 42690 8280 42750 8880
rect 42960 8280 43020 8880
rect 43110 8280 43170 8880
rect 43470 8280 43530 8880
rect 43620 8280 43680 8880
rect 43890 8280 43950 8880
rect 45330 8280 45390 8880
rect 45600 8280 45660 8880
rect 45750 8280 45810 8880
rect 46110 8280 46170 8880
rect 46260 8280 46320 8880
rect 46530 8280 46590 8880
rect 47820 8280 47880 8880
rect 47970 8280 48030 8880
rect 49260 8280 49320 8880
rect 49410 8280 49470 8880
rect 5730 7320 5790 7920
rect 6000 7320 6060 7920
rect 6150 7320 6210 7920
rect 6510 7320 6570 7920
rect 6660 7320 6720 7920
rect 6930 7320 6990 7920
rect 8130 7620 8190 7920
rect 8850 7320 8910 7920
rect 9090 7320 9150 7920
rect 9330 7320 9390 7920
rect 10050 7320 10110 7920
rect 10200 7320 10260 7920
rect 11010 7320 11070 7920
rect 11250 7320 11310 7920
rect 11490 7320 11550 7920
rect 12450 7320 12510 7920
rect 12600 7320 12660 7920
rect 13980 7320 14040 7920
rect 14130 7320 14190 7920
rect 14370 7620 14430 7920
rect 15570 7620 15630 7920
rect 15810 7620 15870 7920
rect 18210 7620 18270 7920
rect 18450 7620 18510 7920
rect 20850 7320 20910 7920
rect 21000 7320 21060 7920
rect 23490 7320 23550 7920
rect 23640 7320 23700 7920
rect 25890 7320 25950 7920
rect 26160 7320 26220 7920
rect 26310 7320 26370 7920
rect 26670 7320 26730 7920
rect 26820 7320 26880 7920
rect 27090 7320 27150 7920
rect 28050 7320 28110 7920
rect 28200 7320 28260 7920
rect 29250 7320 29310 7920
rect 29400 7320 29460 7920
rect 30210 7320 30270 7920
rect 30480 7320 30540 7920
rect 30630 7320 30690 7920
rect 30990 7320 31050 7920
rect 31140 7320 31200 7920
rect 31410 7320 31470 7920
rect 32130 7320 32190 7920
rect 32370 7320 32430 7920
rect 32610 7320 32670 7920
rect 33330 7320 33390 7920
rect 33480 7320 33540 7920
rect 34860 7320 34920 7920
rect 35010 7320 35070 7920
rect 36210 7320 36270 7920
rect 36360 7320 36420 7920
rect 37650 7320 37710 7920
rect 37890 7320 37950 7920
rect 38130 7320 38190 7920
rect 39090 7320 39150 7920
rect 39240 7320 39300 7920
rect 40530 7320 40590 7920
rect 40680 7320 40740 7920
rect 43410 7620 43470 7920
rect 43650 7620 43710 7920
rect 44670 7320 44730 7920
rect 44820 7320 44880 7920
rect 45180 7320 45240 7920
rect 45330 7320 45390 7920
rect 46530 7620 46590 7920
rect 47490 7320 47550 7920
rect 47730 7320 47790 7920
rect 47970 7320 48030 7920
<< ptransistor >>
rect 5820 41280 5880 41880
rect 6060 41280 6120 42480
rect 6210 41280 6270 42480
rect 6930 41280 6990 41880
rect 7170 41280 7230 41880
rect 7980 41280 8040 41880
rect 8220 41280 8280 42480
rect 8370 41280 8430 42480
rect 9090 41280 9150 42480
rect 9360 41280 9420 42480
rect 9510 41280 9570 42480
rect 9870 41280 9930 42480
rect 10020 41280 10080 42480
rect 10290 41280 10350 42480
rect 11100 41280 11160 42480
rect 11250 41280 11310 42480
rect 12540 41280 12600 42480
rect 12690 41280 12750 42480
rect 13890 41280 13950 42480
rect 14040 41280 14100 42480
rect 14280 41280 14340 41880
rect 15570 41280 15630 41880
rect 15810 41280 15870 41880
rect 17250 41280 17310 42480
rect 17400 41280 17460 42480
rect 17640 41280 17700 41880
rect 19410 41280 19470 42480
rect 19680 41280 19740 42480
rect 19830 41280 19890 42480
rect 20190 41280 20250 42480
rect 20340 41280 20400 42480
rect 20610 41280 20670 42480
rect 21330 41280 21390 41880
rect 22770 41280 22830 42480
rect 23040 41280 23100 42480
rect 23190 41280 23250 42480
rect 23550 41280 23610 42480
rect 23700 41280 23760 42480
rect 23970 41280 24030 42480
rect 25260 41280 25320 41880
rect 25500 41280 25560 42480
rect 25650 41280 25710 42480
rect 26850 41280 26910 41880
rect 27090 41280 27150 41880
rect 28050 41280 28110 42480
rect 28200 41280 28260 42480
rect 28440 41280 28500 41880
rect 29250 41280 29310 41880
rect 29490 41280 29550 41880
rect 30450 41280 30510 42480
rect 30600 41280 30660 42480
rect 30840 41280 30900 41880
rect 31890 41280 31950 42480
rect 32040 41280 32100 42480
rect 32280 41280 32340 41880
rect 33330 41280 33390 41880
rect 33570 41280 33630 41880
rect 34770 41280 34830 42480
rect 34920 41280 34980 42480
rect 35970 41280 36030 42480
rect 36240 41280 36300 42480
rect 36390 41280 36450 42480
rect 36750 41280 36810 42480
rect 36900 41280 36960 42480
rect 37170 41280 37230 42480
rect 37980 41280 38040 41880
rect 38220 41280 38280 42480
rect 38370 41280 38430 42480
rect 39570 41280 39630 42480
rect 39840 41280 39900 42480
rect 39990 41280 40050 42480
rect 40350 41280 40410 42480
rect 40500 41280 40560 42480
rect 40770 41280 40830 42480
rect 41970 41280 42030 41880
rect 43170 41280 43230 42480
rect 43320 41280 43380 42480
rect 43560 41280 43620 41880
rect 44370 41280 44430 42480
rect 44520 41280 44580 42480
rect 44760 41280 44820 41880
rect 45330 41280 45390 41880
rect 45810 41280 45870 42480
rect 46080 41280 46140 42480
rect 46230 41280 46290 42480
rect 46590 41280 46650 42480
rect 46740 41280 46800 42480
rect 47010 41280 47070 42480
rect 47490 41280 47550 42480
rect 47760 41280 47820 42480
rect 47910 41280 47970 42480
rect 48270 41280 48330 42480
rect 48420 41280 48480 42480
rect 48690 41280 48750 42480
rect 5970 39720 6030 40920
rect 6210 39720 6270 40920
rect 6450 39720 6510 40920
rect 8370 40320 8430 40920
rect 8610 40320 8670 40920
rect 9810 40320 9870 40920
rect 10050 40320 10110 40920
rect 10770 39720 10830 40920
rect 11010 39720 11070 40920
rect 11250 39720 11310 40920
rect 11730 39720 11790 40920
rect 12000 39720 12060 40920
rect 12150 39720 12210 40920
rect 12510 39720 12570 40920
rect 12660 39720 12720 40920
rect 12930 39720 12990 40920
rect 13650 40320 13710 40920
rect 13890 40320 13950 40920
rect 14610 40320 14670 40920
rect 14850 40320 14910 40920
rect 15090 40320 15150 40920
rect 15810 40320 15870 40920
rect 16530 39720 16590 40920
rect 16680 39720 16740 40920
rect 16920 40320 16980 40920
rect 17820 40320 17880 40920
rect 18060 39720 18120 40920
rect 18210 39720 18270 40920
rect 18690 40320 18750 40920
rect 19410 39720 19470 40920
rect 19560 39720 19620 40920
rect 19800 40320 19860 40920
rect 21090 40320 21150 40920
rect 21330 40320 21390 40920
rect 22050 39720 22110 40920
rect 22320 39720 22380 40920
rect 22470 39720 22530 40920
rect 22830 39720 22890 40920
rect 22980 39720 23040 40920
rect 23250 39720 23310 40920
rect 23970 39720 24030 40920
rect 24120 39720 24180 40920
rect 24930 39720 24990 40920
rect 25080 39720 25140 40920
rect 25320 40320 25380 40920
rect 26370 39720 26430 40920
rect 26610 39720 26670 40920
rect 26850 39720 26910 40920
rect 27090 39720 27150 40920
rect 28050 40320 28110 40920
rect 30690 40320 30750 40920
rect 30930 40320 30990 40920
rect 32130 40320 32190 40920
rect 32370 40320 32430 40920
rect 33570 39720 33630 40920
rect 33840 39720 33900 40920
rect 33990 39720 34050 40920
rect 34350 39720 34410 40920
rect 34500 39720 34560 40920
rect 34770 39720 34830 40920
rect 36210 39720 36270 40920
rect 36360 39720 36420 40920
rect 36600 40320 36660 40920
rect 37890 40320 37950 40920
rect 38130 40320 38190 40920
rect 39090 39720 39150 40920
rect 39240 39720 39300 40920
rect 39480 40320 39540 40920
rect 40530 40320 40590 40920
rect 40770 40320 40830 40920
rect 41970 40320 42030 40920
rect 43170 39720 43230 40920
rect 43320 39720 43380 40920
rect 43560 40320 43620 40920
rect 44850 40320 44910 40920
rect 46140 40320 46200 40920
rect 46380 39720 46440 40920
rect 46530 39720 46590 40920
rect 47730 39720 47790 40920
rect 47880 39720 47940 40920
rect 48120 40320 48180 40920
rect 49410 40320 49470 40920
rect 49650 40320 49710 40920
rect 5730 35280 5790 35880
rect 5970 35280 6030 35880
rect 7170 35280 7230 35880
rect 8460 35280 8520 35880
rect 8700 35280 8760 36480
rect 8850 35280 8910 36480
rect 11010 35280 11070 35880
rect 11250 35280 11310 35880
rect 12300 35280 12360 35880
rect 12540 35280 12600 36480
rect 12690 35280 12750 36480
rect 15180 35280 15240 35880
rect 15420 35280 15480 36480
rect 15570 35280 15630 36480
rect 16770 35280 16830 35880
rect 17010 35280 17070 35880
rect 17250 35280 17310 35880
rect 18210 35280 18270 35880
rect 18450 35280 18510 35880
rect 19650 35280 19710 35880
rect 19890 35280 19950 35880
rect 21090 35280 21150 35880
rect 21330 35280 21390 35880
rect 22530 35280 22590 35880
rect 22770 35280 22830 35880
rect 23970 35280 24030 35880
rect 25170 35280 25230 35880
rect 25410 35280 25470 35880
rect 26610 35280 26670 36480
rect 26760 35280 26820 36480
rect 27000 35280 27060 35880
rect 28050 35280 28110 35880
rect 28290 35280 28350 35880
rect 29250 35280 29310 35880
rect 29490 35280 29550 35880
rect 30210 35280 30270 36480
rect 30360 35280 30420 36480
rect 30600 35280 30660 35880
rect 31410 35280 31470 35880
rect 32220 35280 32280 35880
rect 32460 35280 32520 36480
rect 32610 35280 32670 36480
rect 33330 35280 33390 35880
rect 33570 35280 33630 35880
rect 34770 35280 34830 35880
rect 35010 35280 35070 35880
rect 35730 35280 35790 36480
rect 36000 35280 36060 36480
rect 36150 35280 36210 36480
rect 36510 35280 36570 36480
rect 36660 35280 36720 36480
rect 36930 35280 36990 36480
rect 39090 35280 39150 35880
rect 40050 35280 40110 36480
rect 40290 35280 40350 36480
rect 40530 35280 40590 36480
rect 40770 35280 40830 36480
rect 41730 35280 41790 35880
rect 42540 35280 42600 35880
rect 42780 35280 42840 36480
rect 42930 35280 42990 36480
rect 43650 35280 43710 35880
rect 44610 35280 44670 36480
rect 44760 35280 44820 36480
rect 45000 35280 45060 35880
rect 46290 35280 46350 35880
rect 46530 35280 46590 35880
rect 47730 35280 47790 36480
rect 47880 35280 47940 36480
rect 48120 35280 48180 35880
rect 49410 35280 49470 35880
rect 49650 35280 49710 35880
rect 6780 34320 6840 34920
rect 7020 33720 7080 34920
rect 7170 33720 7230 34920
rect 7980 34320 8040 34920
rect 8220 33720 8280 34920
rect 8370 33720 8430 34920
rect 9090 33720 9150 34920
rect 9360 33720 9420 34920
rect 9510 33720 9570 34920
rect 9870 33720 9930 34920
rect 10020 33720 10080 34920
rect 10290 33720 10350 34920
rect 11250 33720 11310 34920
rect 11520 33720 11580 34920
rect 11670 33720 11730 34920
rect 12030 33720 12090 34920
rect 12180 33720 12240 34920
rect 12450 33720 12510 34920
rect 13890 34320 13950 34920
rect 15330 34320 15390 34920
rect 15570 34320 15630 34920
rect 16770 33720 16830 34920
rect 16920 33720 16980 34920
rect 17160 34320 17220 34920
rect 19410 34320 19470 34920
rect 19650 34320 19710 34920
rect 20850 34320 20910 34920
rect 21090 34320 21150 34920
rect 21330 34320 21390 34920
rect 23490 33720 23550 34920
rect 23640 33720 23700 34920
rect 23880 34320 23940 34920
rect 24930 33720 24990 34920
rect 25080 33720 25140 34920
rect 25320 34320 25380 34920
rect 26130 33720 26190 34920
rect 26400 33720 26460 34920
rect 26550 33720 26610 34920
rect 26910 33720 26970 34920
rect 27060 33720 27120 34920
rect 27330 33720 27390 34920
rect 30450 34320 30510 34920
rect 31170 34320 31230 34920
rect 31410 34320 31470 34920
rect 32130 33720 32190 34920
rect 32280 33720 32340 34920
rect 32520 34320 32580 34920
rect 33330 34320 33390 34920
rect 33570 34320 33630 34920
rect 34770 34320 34830 34920
rect 35010 34320 35070 34920
rect 36210 34320 36270 34920
rect 36450 34320 36510 34920
rect 37650 34320 37710 34920
rect 37890 34320 37950 34920
rect 39090 34320 39150 34920
rect 39330 34320 39390 34920
rect 40290 33720 40350 34920
rect 40440 33720 40500 34920
rect 40680 34320 40740 34920
rect 41730 34320 41790 34920
rect 41970 34320 42030 34920
rect 43170 33720 43230 34920
rect 43320 33720 43380 34920
rect 43560 34320 43620 34920
rect 44370 33720 44430 34920
rect 44640 33720 44700 34920
rect 44790 33720 44850 34920
rect 45150 33720 45210 34920
rect 45300 33720 45360 34920
rect 45570 33720 45630 34920
rect 46290 33720 46350 34920
rect 46440 33720 46500 34920
rect 46680 34320 46740 34920
rect 47730 34320 47790 34920
rect 47970 34320 48030 34920
rect 49170 34320 49230 34920
rect 49410 34320 49470 34920
rect 5490 29280 5550 30480
rect 5760 29280 5820 30480
rect 5910 29280 5970 30480
rect 6270 29280 6330 30480
rect 6420 29280 6480 30480
rect 6690 29280 6750 30480
rect 8130 29280 8190 30480
rect 8280 29280 8340 30480
rect 8520 29280 8580 29880
rect 9810 29280 9870 29880
rect 10050 29280 10110 29880
rect 11250 29280 11310 30480
rect 11520 29280 11580 30480
rect 11670 29280 11730 30480
rect 12030 29280 12090 30480
rect 12180 29280 12240 30480
rect 12450 29280 12510 30480
rect 14850 29280 14910 30480
rect 15120 29280 15180 30480
rect 15270 29280 15330 30480
rect 15630 29280 15690 30480
rect 15780 29280 15840 30480
rect 16050 29280 16110 30480
rect 17250 29280 17310 30480
rect 17520 29280 17580 30480
rect 17670 29280 17730 30480
rect 18030 29280 18090 30480
rect 18180 29280 18240 30480
rect 18450 29280 18510 30480
rect 19410 29280 19470 30480
rect 19680 29280 19740 30480
rect 19830 29280 19890 30480
rect 20190 29280 20250 30480
rect 20340 29280 20400 30480
rect 20610 29280 20670 30480
rect 21330 29280 21390 29880
rect 21570 29280 21630 29880
rect 22380 29280 22440 29880
rect 22620 29280 22680 30480
rect 22770 29280 22830 30480
rect 23970 29280 24030 29880
rect 24930 29280 24990 29880
rect 25170 29280 25230 29880
rect 25410 29280 25470 29880
rect 26220 29280 26280 29880
rect 26460 29280 26520 30480
rect 26610 29280 26670 30480
rect 27330 29280 27390 29880
rect 27810 29280 27870 29880
rect 28050 29280 28110 29880
rect 28770 29280 28830 29880
rect 29340 29280 29400 29880
rect 29580 29280 29640 30480
rect 29730 29280 29790 30480
rect 30930 29280 30990 30480
rect 31200 29280 31260 30480
rect 31350 29280 31410 30480
rect 31710 29280 31770 30480
rect 31860 29280 31920 30480
rect 32130 29280 32190 30480
rect 33330 29280 33390 29880
rect 33570 29280 33630 29880
rect 34770 29280 34830 29880
rect 35010 29280 35070 29880
rect 36300 29280 36360 29880
rect 36540 29280 36600 30480
rect 36690 29280 36750 30480
rect 37890 29280 37950 29880
rect 38130 29280 38190 29880
rect 39090 29280 39150 30480
rect 39240 29280 39300 30480
rect 39480 29280 39540 29880
rect 40770 29280 40830 29880
rect 41730 29280 41790 29880
rect 41970 29280 42030 29880
rect 43260 29280 43320 29880
rect 43500 29280 43560 30480
rect 43650 29280 43710 30480
rect 44610 29280 44670 30480
rect 44760 29280 44820 30480
rect 45000 29280 45060 29880
rect 46290 29280 46350 29880
rect 46530 29280 46590 29880
rect 48210 29280 48270 30480
rect 48480 29280 48540 30480
rect 48630 29280 48690 30480
rect 48990 29280 49050 30480
rect 49140 29280 49200 30480
rect 49410 29280 49470 30480
rect 7170 27720 7230 28920
rect 7440 27720 7500 28920
rect 7590 27720 7650 28920
rect 7950 27720 8010 28920
rect 8100 27720 8160 28920
rect 8370 27720 8430 28920
rect 8850 28320 8910 28920
rect 9090 28320 9150 28920
rect 9570 27720 9630 28920
rect 9840 27720 9900 28920
rect 9990 27720 10050 28920
rect 10350 27720 10410 28920
rect 10500 27720 10560 28920
rect 10770 27720 10830 28920
rect 11250 27720 11310 28920
rect 11400 27720 11460 28920
rect 11640 28320 11700 28920
rect 12210 28320 12270 28920
rect 12450 28320 12510 28920
rect 12930 28320 12990 28920
rect 13170 28320 13230 28920
rect 13890 28320 13950 28920
rect 14130 28320 14190 28920
rect 14370 28320 14430 28920
rect 15570 28320 15630 28920
rect 15810 28320 15870 28920
rect 16770 28320 16830 28920
rect 17010 28320 17070 28920
rect 18210 28320 18270 28920
rect 18450 28320 18510 28920
rect 19500 28320 19560 28920
rect 19740 27720 19800 28920
rect 19890 27720 19950 28920
rect 21090 28320 21150 28920
rect 21330 28320 21390 28920
rect 22290 28320 22350 28920
rect 22530 28320 22590 28920
rect 23730 28320 23790 28920
rect 23970 28320 24030 28920
rect 25170 28320 25230 28920
rect 25410 28320 25470 28920
rect 26610 28320 26670 28920
rect 26850 28320 26910 28920
rect 28620 28320 28680 28920
rect 28860 27720 28920 28920
rect 29010 27720 29070 28920
rect 30450 28320 30510 28920
rect 30690 28320 30750 28920
rect 31980 28320 32040 28920
rect 32220 27720 32280 28920
rect 32370 27720 32430 28920
rect 33090 27720 33150 28920
rect 33360 27720 33420 28920
rect 33510 27720 33570 28920
rect 33870 27720 33930 28920
rect 34020 27720 34080 28920
rect 34290 27720 34350 28920
rect 35010 28320 35070 28920
rect 35250 28320 35310 28920
rect 36210 28320 36270 28920
rect 36450 28320 36510 28920
rect 37650 28320 37710 28920
rect 37890 28320 37950 28920
rect 38850 28320 38910 28920
rect 39090 28320 39150 28920
rect 39810 27720 39870 28920
rect 40080 27720 40140 28920
rect 40230 27720 40290 28920
rect 40590 27720 40650 28920
rect 40740 27720 40800 28920
rect 41010 27720 41070 28920
rect 41730 28320 41790 28920
rect 41970 28320 42030 28920
rect 43260 28320 43320 28920
rect 43500 27720 43560 28920
rect 43650 27720 43710 28920
rect 44610 27720 44670 28920
rect 44760 27720 44820 28920
rect 45000 28320 45060 28920
rect 46050 27720 46110 28920
rect 46200 27720 46260 28920
rect 46440 28320 46500 28920
rect 47010 28320 47070 28920
rect 47490 27720 47550 28920
rect 47730 27720 47790 28920
rect 47970 27720 48030 28920
rect 48210 27720 48270 28920
rect 48690 28320 48750 28920
rect 48930 28320 48990 28920
rect 49410 27720 49470 28920
rect 49560 27720 49620 28920
rect 49800 28320 49860 28920
rect 5490 23280 5550 24480
rect 5760 23280 5820 24480
rect 5910 23280 5970 24480
rect 6270 23280 6330 24480
rect 6420 23280 6480 24480
rect 6690 23280 6750 24480
rect 7170 23280 7230 23880
rect 7410 23280 7470 23880
rect 7980 23280 8040 23880
rect 8220 23280 8280 24480
rect 8370 23280 8430 24480
rect 8850 23280 8910 23880
rect 9090 23280 9150 23880
rect 9570 23280 9630 24480
rect 9840 23280 9900 24480
rect 9990 23280 10050 24480
rect 10350 23280 10410 24480
rect 10500 23280 10560 24480
rect 10770 23280 10830 24480
rect 12210 23280 12270 24480
rect 12450 23280 12510 24480
rect 12690 23280 12750 24480
rect 13890 23280 13950 23880
rect 15180 23280 15240 23880
rect 15420 23280 15480 24480
rect 15570 23280 15630 24480
rect 20850 23280 20910 23880
rect 21090 23280 21150 23880
rect 23250 23280 23310 23880
rect 23490 23280 23550 23880
rect 25650 23280 25710 24480
rect 25920 23280 25980 24480
rect 26070 23280 26130 24480
rect 26430 23280 26490 24480
rect 26580 23280 26640 24480
rect 26850 23280 26910 24480
rect 28140 23280 28200 23880
rect 28380 23280 28440 24480
rect 28530 23280 28590 24480
rect 30450 23280 30510 23880
rect 31260 23280 31320 23880
rect 31500 23280 31560 24480
rect 31650 23280 31710 24480
rect 32370 23280 32430 23880
rect 33330 23280 33390 23880
rect 33570 23280 33630 23880
rect 34770 23280 34830 23880
rect 35010 23280 35070 23880
rect 36210 23280 36270 23880
rect 36450 23280 36510 23880
rect 37650 23280 37710 23880
rect 37890 23280 37950 23880
rect 39090 23280 39150 23880
rect 39330 23280 39390 23880
rect 40530 23280 40590 23880
rect 40770 23280 40830 23880
rect 41970 23280 42030 23880
rect 42210 23280 42270 23880
rect 43410 23280 43470 24480
rect 43560 23280 43620 24480
rect 44610 23280 44670 23880
rect 47970 23280 48030 24480
rect 48240 23280 48300 24480
rect 48390 23280 48450 24480
rect 48750 23280 48810 24480
rect 48900 23280 48960 24480
rect 49170 23280 49230 24480
rect 5490 21720 5550 22920
rect 5760 21720 5820 22920
rect 5910 21720 5970 22920
rect 6270 21720 6330 22920
rect 6420 21720 6480 22920
rect 6690 21720 6750 22920
rect 8370 22320 8430 22920
rect 8610 22320 8670 22920
rect 9810 22320 9870 22920
rect 10050 22320 10110 22920
rect 11340 22320 11400 22920
rect 11580 21720 11640 22920
rect 11730 21720 11790 22920
rect 14370 21720 14430 22920
rect 14640 21720 14700 22920
rect 14790 21720 14850 22920
rect 15150 21720 15210 22920
rect 15300 21720 15360 22920
rect 15570 21720 15630 22920
rect 17010 22320 17070 22920
rect 18210 22320 18270 22920
rect 18450 22320 18510 22920
rect 18930 21720 18990 22920
rect 19200 21720 19260 22920
rect 19350 21720 19410 22920
rect 19710 21720 19770 22920
rect 19860 21720 19920 22920
rect 20130 21720 20190 22920
rect 20610 21720 20670 22920
rect 20880 21720 20940 22920
rect 21030 21720 21090 22920
rect 21390 21720 21450 22920
rect 21540 21720 21600 22920
rect 21810 21720 21870 22920
rect 22380 22320 22440 22920
rect 22620 21720 22680 22920
rect 22770 21720 22830 22920
rect 25170 22320 25230 22920
rect 26460 22320 26520 22920
rect 26700 21720 26760 22920
rect 26850 21720 26910 22920
rect 28140 22320 28200 22920
rect 28380 21720 28440 22920
rect 28530 21720 28590 22920
rect 29250 22320 29310 22920
rect 29490 22320 29550 22920
rect 30450 21720 30510 22920
rect 30600 21720 30660 22920
rect 30840 22320 30900 22920
rect 32130 22320 32190 22920
rect 32370 22320 32430 22920
rect 33330 22320 33390 22920
rect 33570 22320 33630 22920
rect 34770 22320 34830 22920
rect 35010 22320 35070 22920
rect 35970 22320 36030 22920
rect 36210 22320 36270 22920
rect 36930 21720 36990 22920
rect 37200 21720 37260 22920
rect 37350 21720 37410 22920
rect 37710 21720 37770 22920
rect 37860 21720 37920 22920
rect 38130 21720 38190 22920
rect 39180 22320 39240 22920
rect 39420 21720 39480 22920
rect 39570 21720 39630 22920
rect 40530 22320 40590 22920
rect 40770 22320 40830 22920
rect 41820 22320 41880 22920
rect 42060 21720 42120 22920
rect 42210 21720 42270 22920
rect 43410 21720 43470 22920
rect 43560 21720 43620 22920
rect 44370 21720 44430 22920
rect 44640 21720 44700 22920
rect 44790 21720 44850 22920
rect 45150 21720 45210 22920
rect 45300 21720 45360 22920
rect 45570 21720 45630 22920
rect 46050 21720 46110 22920
rect 46320 21720 46380 22920
rect 46470 21720 46530 22920
rect 46830 21720 46890 22920
rect 46980 21720 47040 22920
rect 47250 21720 47310 22920
rect 47730 22320 47790 22920
rect 48930 21720 48990 22920
rect 49170 21720 49230 22920
rect 49410 21720 49470 22920
rect 49650 21720 49710 22920
rect 5820 17280 5880 17880
rect 6060 17280 6120 18480
rect 6210 17280 6270 18480
rect 9090 17280 9150 18480
rect 9360 17280 9420 18480
rect 9510 17280 9570 18480
rect 9870 17280 9930 18480
rect 10020 17280 10080 18480
rect 10290 17280 10350 18480
rect 11730 17280 11790 18480
rect 12000 17280 12060 18480
rect 12150 17280 12210 18480
rect 12510 17280 12570 18480
rect 12660 17280 12720 18480
rect 12930 17280 12990 18480
rect 13650 17280 13710 18480
rect 13920 17280 13980 18480
rect 14070 17280 14130 18480
rect 14430 17280 14490 18480
rect 14580 17280 14640 18480
rect 14850 17280 14910 18480
rect 15570 17280 15630 18480
rect 15810 17280 15870 18480
rect 16050 17280 16110 18480
rect 18060 17280 18120 17880
rect 18300 17280 18360 18480
rect 18450 17280 18510 18480
rect 19650 17280 19710 17880
rect 19890 17280 19950 17880
rect 21090 17280 21150 17880
rect 21330 17280 21390 17880
rect 22290 17280 22350 17880
rect 22530 17280 22590 17880
rect 23730 17280 23790 17880
rect 23970 17280 24030 17880
rect 24690 17280 24750 18480
rect 24960 17280 25020 18480
rect 25110 17280 25170 18480
rect 25470 17280 25530 18480
rect 25620 17280 25680 18480
rect 25890 17280 25950 18480
rect 26370 17280 26430 18480
rect 26520 17280 26580 18480
rect 26760 17280 26820 17880
rect 27330 17280 27390 17880
rect 28620 17280 28680 17880
rect 28860 17280 28920 18480
rect 29010 17280 29070 18480
rect 30690 17280 30750 17880
rect 30930 17280 30990 17880
rect 32130 17280 32190 17880
rect 32370 17280 32430 17880
rect 33330 17280 33390 18480
rect 33480 17280 33540 18480
rect 33720 17280 33780 17880
rect 35970 17280 36030 17880
rect 36210 17280 36270 17880
rect 36930 17280 36990 18480
rect 37170 17280 37230 18480
rect 37410 17280 37470 18480
rect 38130 17280 38190 17880
rect 38370 17280 38430 17880
rect 39090 17280 39150 17880
rect 39330 17280 39390 17880
rect 40530 17280 40590 17880
rect 40770 17280 40830 17880
rect 41730 17280 41790 17880
rect 42930 17280 42990 18480
rect 43170 17280 43230 18480
rect 43410 17280 43470 18480
rect 43650 17280 43710 18480
rect 44610 17280 44670 18480
rect 44760 17280 44820 18480
rect 45000 17280 45060 17880
rect 46290 17280 46350 17880
rect 46530 17280 46590 17880
rect 47730 17280 47790 18480
rect 47880 17280 47940 18480
rect 49170 17280 49230 18480
rect 49320 17280 49380 18480
rect 49560 17280 49620 17880
rect 6450 16320 6510 16920
rect 6690 16320 6750 16920
rect 7890 15720 7950 16920
rect 8160 15720 8220 16920
rect 8310 15720 8370 16920
rect 8670 15720 8730 16920
rect 8820 15720 8880 16920
rect 9090 15720 9150 16920
rect 9570 15720 9630 16920
rect 9840 15720 9900 16920
rect 9990 15720 10050 16920
rect 10350 15720 10410 16920
rect 10500 15720 10560 16920
rect 10770 15720 10830 16920
rect 11250 15720 11310 16920
rect 11520 15720 11580 16920
rect 11670 15720 11730 16920
rect 12030 15720 12090 16920
rect 12180 15720 12240 16920
rect 12450 15720 12510 16920
rect 13410 15720 13470 16920
rect 13680 15720 13740 16920
rect 13830 15720 13890 16920
rect 14190 15720 14250 16920
rect 14340 15720 14400 16920
rect 14610 15720 14670 16920
rect 15090 15720 15150 16920
rect 15360 15720 15420 16920
rect 15510 15720 15570 16920
rect 15870 15720 15930 16920
rect 16020 15720 16080 16920
rect 16290 15720 16350 16920
rect 16770 15720 16830 16920
rect 17010 15720 17070 16920
rect 17250 15720 17310 16920
rect 17730 16320 17790 16920
rect 18300 16320 18360 16920
rect 18540 15720 18600 16920
rect 18690 15720 18750 16920
rect 19410 16320 19470 16920
rect 19650 16320 19710 16920
rect 20850 15720 20910 16920
rect 21000 15720 21060 16920
rect 21240 16320 21300 16920
rect 22380 16320 22440 16920
rect 22620 15720 22680 16920
rect 22770 15720 22830 16920
rect 23730 16320 23790 16920
rect 23970 16320 24030 16920
rect 24930 16320 24990 16920
rect 25170 16320 25230 16920
rect 25890 15720 25950 16920
rect 26160 15720 26220 16920
rect 26310 15720 26370 16920
rect 26670 15720 26730 16920
rect 26820 15720 26880 16920
rect 27090 15720 27150 16920
rect 28050 16320 28110 16920
rect 28290 16320 28350 16920
rect 29250 16320 29310 16920
rect 29490 16320 29550 16920
rect 30450 15720 30510 16920
rect 30720 15720 30780 16920
rect 30870 15720 30930 16920
rect 31230 15720 31290 16920
rect 31380 15720 31440 16920
rect 31650 15720 31710 16920
rect 32370 16320 32430 16920
rect 32610 16320 32670 16920
rect 33330 16320 33390 16920
rect 33570 16320 33630 16920
rect 34770 16320 34830 16920
rect 35010 16320 35070 16920
rect 36210 15720 36270 16920
rect 36360 15720 36420 16920
rect 36600 16320 36660 16920
rect 37890 16320 37950 16920
rect 38130 16320 38190 16920
rect 38850 15720 38910 16920
rect 39120 15720 39180 16920
rect 39270 15720 39330 16920
rect 39630 15720 39690 16920
rect 39780 15720 39840 16920
rect 40050 15720 40110 16920
rect 41730 15720 41790 16920
rect 42000 15720 42060 16920
rect 42150 15720 42210 16920
rect 42510 15720 42570 16920
rect 42660 15720 42720 16920
rect 42930 15720 42990 16920
rect 44610 15720 44670 16920
rect 44760 15720 44820 16920
rect 45000 16320 45060 16920
rect 46290 16320 46350 16920
rect 46530 16320 46590 16920
rect 47730 16320 47790 16920
rect 47970 16320 48030 16920
rect 49170 15720 49230 16920
rect 49320 15720 49380 16920
rect 49560 16320 49620 16920
rect 6930 11280 6990 11880
rect 7170 11280 7230 11880
rect 9090 11280 9150 12480
rect 9240 11280 9300 12480
rect 9660 11280 9720 12480
rect 9810 11280 9870 12480
rect 11010 11280 11070 11880
rect 11250 11280 11310 11880
rect 12300 11280 12360 11880
rect 12540 11280 12600 12480
rect 12690 11280 12750 12480
rect 16050 11280 16110 11880
rect 16290 11280 16350 11880
rect 16860 11280 16920 11880
rect 17100 11280 17160 12480
rect 17250 11280 17310 12480
rect 17730 11280 17790 12480
rect 18000 11280 18060 12480
rect 18150 11280 18210 12480
rect 18510 11280 18570 12480
rect 18660 11280 18720 12480
rect 18930 11280 18990 12480
rect 19410 11280 19470 12480
rect 19680 11280 19740 12480
rect 19830 11280 19890 12480
rect 20190 11280 20250 12480
rect 20340 11280 20400 12480
rect 20610 11280 20670 12480
rect 22050 11280 22110 12480
rect 22320 11280 22380 12480
rect 22470 11280 22530 12480
rect 22830 11280 22890 12480
rect 22980 11280 23040 12480
rect 23250 11280 23310 12480
rect 25170 11280 25230 12480
rect 25320 11280 25380 12480
rect 25560 11280 25620 11880
rect 26850 11280 26910 11880
rect 27090 11280 27150 11880
rect 29250 11280 29310 12480
rect 29400 11280 29460 12480
rect 29640 11280 29700 11880
rect 30540 11280 30600 11880
rect 30780 11280 30840 12480
rect 30930 11280 30990 12480
rect 32130 11280 32190 11880
rect 32370 11280 32430 11880
rect 33090 11280 33150 12480
rect 33360 11280 33420 12480
rect 33510 11280 33570 12480
rect 33870 11280 33930 12480
rect 34020 11280 34080 12480
rect 34290 11280 34350 12480
rect 34770 11280 34830 12480
rect 34920 11280 34980 12480
rect 35160 11280 35220 11880
rect 36210 11280 36270 11880
rect 36450 11280 36510 11880
rect 37650 11280 37710 11880
rect 37890 11280 37950 11880
rect 39090 11280 39150 11880
rect 39330 11280 39390 11880
rect 40380 11280 40440 11880
rect 40620 11280 40680 12480
rect 40770 11280 40830 12480
rect 41730 11280 41790 11880
rect 41970 11280 42030 11880
rect 42210 11280 42270 11880
rect 43410 11280 43470 11880
rect 43650 11280 43710 11880
rect 44610 11280 44670 12480
rect 44760 11280 44820 12480
rect 45000 11280 45060 11880
rect 46290 11280 46350 11880
rect 46530 11280 46590 11880
rect 47730 11280 47790 12480
rect 47880 11280 47940 12480
rect 48120 11280 48180 11880
rect 49410 11280 49470 11880
rect 49650 11280 49710 11880
rect 5820 10320 5880 10920
rect 6060 9720 6120 10920
rect 6210 9720 6270 10920
rect 6930 10320 6990 10920
rect 7170 10320 7230 10920
rect 7890 9720 7950 10920
rect 8160 9720 8220 10920
rect 8310 9720 8370 10920
rect 8670 9720 8730 10920
rect 8820 9720 8880 10920
rect 9090 9720 9150 10920
rect 9810 10320 9870 10920
rect 10050 10320 10110 10920
rect 10290 10320 10350 10920
rect 11490 10320 11550 10920
rect 11730 10320 11790 10920
rect 13890 9720 13950 10920
rect 14160 9720 14220 10920
rect 14310 9720 14370 10920
rect 14670 9720 14730 10920
rect 14820 9720 14880 10920
rect 15090 9720 15150 10920
rect 16530 10320 16590 10920
rect 16770 10320 16830 10920
rect 17490 9720 17550 10920
rect 17760 9720 17820 10920
rect 17910 9720 17970 10920
rect 18270 9720 18330 10920
rect 18420 9720 18480 10920
rect 18690 9720 18750 10920
rect 19410 9720 19470 10920
rect 19680 9720 19740 10920
rect 19830 9720 19890 10920
rect 20190 9720 20250 10920
rect 20340 9720 20400 10920
rect 20610 9720 20670 10920
rect 21330 10320 21390 10920
rect 21570 10320 21630 10920
rect 22050 9720 22110 10920
rect 22320 9720 22380 10920
rect 22470 9720 22530 10920
rect 22830 9720 22890 10920
rect 22980 9720 23040 10920
rect 23250 9720 23310 10920
rect 23970 10320 24030 10920
rect 24210 10320 24270 10920
rect 25650 9720 25710 10920
rect 25920 9720 25980 10920
rect 26070 9720 26130 10920
rect 26430 9720 26490 10920
rect 26580 9720 26640 10920
rect 26850 9720 26910 10920
rect 28050 10320 28110 10920
rect 28290 10320 28350 10920
rect 29490 10320 29550 10920
rect 30690 10320 30750 10920
rect 31890 9720 31950 10920
rect 32040 9720 32100 10920
rect 32280 10320 32340 10920
rect 33330 9720 33390 10920
rect 33600 9720 33660 10920
rect 33750 9720 33810 10920
rect 34110 9720 34170 10920
rect 34260 9720 34320 10920
rect 34530 9720 34590 10920
rect 35730 10320 35790 10920
rect 35970 10320 36030 10920
rect 36210 10320 36270 10920
rect 36930 10320 36990 10920
rect 37170 10320 37230 10920
rect 37890 10320 37950 10920
rect 38130 10320 38190 10920
rect 38370 10320 38430 10920
rect 39090 9720 39150 10920
rect 39240 9720 39300 10920
rect 39480 10320 39540 10920
rect 40530 10320 40590 10920
rect 40770 10320 40830 10920
rect 41730 10320 41790 10920
rect 41970 10320 42030 10920
rect 42690 9720 42750 10920
rect 42960 9720 43020 10920
rect 43110 9720 43170 10920
rect 43470 9720 43530 10920
rect 43620 9720 43680 10920
rect 43890 9720 43950 10920
rect 45330 9720 45390 10920
rect 45600 9720 45660 10920
rect 45750 9720 45810 10920
rect 46110 9720 46170 10920
rect 46260 9720 46320 10920
rect 46530 9720 46590 10920
rect 47730 10320 47790 10920
rect 47970 10320 48030 10920
rect 49170 10320 49230 10920
rect 49410 10320 49470 10920
rect 5730 5280 5790 6480
rect 6000 5280 6060 6480
rect 6150 5280 6210 6480
rect 6510 5280 6570 6480
rect 6660 5280 6720 6480
rect 6930 5280 6990 6480
rect 8130 5280 8190 5880
rect 8940 5280 9000 5880
rect 9180 5280 9240 6480
rect 9330 5280 9390 6480
rect 10050 5280 10110 5880
rect 10290 5280 10350 5880
rect 11100 5280 11160 5880
rect 11340 5280 11400 6480
rect 11490 5280 11550 6480
rect 12450 5280 12510 5880
rect 12690 5280 12750 5880
rect 13890 5280 13950 6480
rect 14130 5280 14190 6480
rect 14370 5280 14430 6480
rect 15570 5280 15630 6480
rect 15720 5280 15780 6480
rect 18210 5280 18270 6480
rect 18360 5280 18420 6480
rect 20850 5280 20910 5880
rect 21090 5280 21150 5880
rect 23490 5280 23550 5880
rect 23730 5280 23790 5880
rect 25890 5280 25950 6480
rect 26160 5280 26220 6480
rect 26310 5280 26370 6480
rect 26670 5280 26730 6480
rect 26820 5280 26880 6480
rect 27090 5280 27150 6480
rect 28050 5280 28110 5880
rect 28290 5280 28350 5880
rect 29250 5280 29310 5880
rect 29490 5280 29550 5880
rect 30210 5280 30270 6480
rect 30480 5280 30540 6480
rect 30630 5280 30690 6480
rect 30990 5280 31050 6480
rect 31140 5280 31200 6480
rect 31410 5280 31470 6480
rect 32130 5280 32190 6480
rect 32280 5280 32340 6480
rect 32520 5280 32580 5880
rect 33330 5280 33390 5880
rect 33570 5280 33630 5880
rect 34770 5280 34830 5880
rect 35010 5280 35070 5880
rect 36210 5280 36270 5880
rect 36450 5280 36510 5880
rect 37740 5280 37800 5880
rect 37980 5280 38040 6480
rect 38130 5280 38190 6480
rect 39090 5280 39150 5880
rect 39330 5280 39390 5880
rect 40530 5280 40590 5880
rect 40770 5280 40830 5880
rect 43410 5280 43470 6480
rect 43560 5280 43620 6480
rect 44610 5280 44670 6480
rect 44850 5280 44910 6480
rect 45090 5280 45150 6480
rect 45330 5280 45390 6480
rect 46530 5280 46590 5880
rect 47580 5280 47640 5880
rect 47820 5280 47880 6480
rect 47970 5280 48030 6480
<< ndiffusion >>
rect 5700 43320 5730 43920
rect 5790 43320 5820 43920
rect 5940 43320 5970 43920
rect 6030 43890 6210 43920
rect 6030 43470 6060 43890
rect 6180 43470 6210 43890
rect 6030 43320 6210 43470
rect 6270 43320 6300 43920
rect 6900 43320 6930 43920
rect 6990 43320 7080 43920
rect 7140 43320 7170 43920
rect 7860 43320 7890 43920
rect 7950 43320 7980 43920
rect 8100 43320 8130 43920
rect 8190 43890 8370 43920
rect 8190 43470 8220 43890
rect 8340 43470 8370 43890
rect 8190 43320 8370 43470
rect 8430 43320 8460 43920
rect 9060 43320 9090 43920
rect 9150 43890 9360 43920
rect 9150 43440 9180 43890
rect 9330 43440 9360 43890
rect 9150 43320 9360 43440
rect 9420 43320 9510 43920
rect 9570 43860 9870 43920
rect 9570 43440 9660 43860
rect 9780 43440 9870 43860
rect 9570 43320 9870 43440
rect 9930 43320 10020 43920
rect 10080 43890 10290 43920
rect 10080 43440 10110 43890
rect 10260 43440 10290 43890
rect 10080 43320 10290 43440
rect 10350 43320 10380 43920
rect 10980 43620 11010 43920
rect 11070 43620 11100 43920
rect 11220 43620 11250 43920
rect 11310 43620 11340 43920
rect 12420 43620 12450 43920
rect 12510 43620 12540 43920
rect 12660 43620 12690 43920
rect 12750 43620 12780 43920
rect 13860 43320 13890 43920
rect 13950 43890 14130 43920
rect 13950 43470 13980 43890
rect 14100 43470 14130 43890
rect 13950 43320 14130 43470
rect 14190 43320 14220 43920
rect 14340 43320 14370 43920
rect 14430 43320 14460 43920
rect 15540 43320 15570 43920
rect 15630 43320 15720 43920
rect 15780 43320 15810 43920
rect 17220 43320 17250 43920
rect 17310 43890 17490 43920
rect 17310 43470 17340 43890
rect 17460 43470 17490 43890
rect 17310 43320 17490 43470
rect 17550 43320 17580 43920
rect 17700 43320 17730 43920
rect 17790 43320 17820 43920
rect 19380 43320 19410 43920
rect 19470 43890 19680 43920
rect 19470 43440 19500 43890
rect 19650 43440 19680 43890
rect 19470 43320 19680 43440
rect 19740 43320 19830 43920
rect 19890 43860 20190 43920
rect 19890 43440 19980 43860
rect 20100 43440 20190 43860
rect 19890 43320 20190 43440
rect 20250 43320 20340 43920
rect 20400 43890 20610 43920
rect 20400 43440 20430 43890
rect 20580 43440 20610 43890
rect 20400 43320 20610 43440
rect 20670 43320 20700 43920
rect 21300 43650 21330 43920
rect 21180 43620 21330 43650
rect 21390 43650 21420 43920
rect 21390 43620 21540 43650
rect 22740 43320 22770 43920
rect 22830 43890 23040 43920
rect 22830 43440 22860 43890
rect 23010 43440 23040 43890
rect 22830 43320 23040 43440
rect 23100 43320 23190 43920
rect 23250 43860 23550 43920
rect 23250 43440 23340 43860
rect 23460 43440 23550 43860
rect 23250 43320 23550 43440
rect 23610 43320 23700 43920
rect 23760 43890 23970 43920
rect 23760 43440 23790 43890
rect 23940 43440 23970 43890
rect 23760 43320 23970 43440
rect 24030 43320 24060 43920
rect 25140 43320 25170 43920
rect 25230 43320 25260 43920
rect 25380 43320 25410 43920
rect 25470 43890 25650 43920
rect 25470 43470 25500 43890
rect 25620 43470 25650 43890
rect 25470 43320 25650 43470
rect 25710 43320 25740 43920
rect 26820 43320 26850 43920
rect 26910 43320 27000 43920
rect 27060 43320 27090 43920
rect 28020 43320 28050 43920
rect 28110 43890 28290 43920
rect 28110 43470 28140 43890
rect 28260 43470 28290 43890
rect 28110 43320 28290 43470
rect 28350 43320 28380 43920
rect 28500 43320 28530 43920
rect 28590 43320 28620 43920
rect 29220 43320 29250 43920
rect 29310 43320 29400 43920
rect 29460 43320 29490 43920
rect 30420 43320 30450 43920
rect 30510 43890 30690 43920
rect 30510 43470 30540 43890
rect 30660 43470 30690 43890
rect 30510 43320 30690 43470
rect 30750 43320 30780 43920
rect 30900 43320 30930 43920
rect 30990 43320 31020 43920
rect 31860 43320 31890 43920
rect 31950 43890 32130 43920
rect 31950 43470 31980 43890
rect 32100 43470 32130 43890
rect 31950 43320 32130 43470
rect 32190 43320 32220 43920
rect 32340 43320 32370 43920
rect 32430 43320 32460 43920
rect 33390 43320 33420 43920
rect 33480 43320 33570 43920
rect 33630 43320 33660 43920
rect 34740 43620 34770 43920
rect 34830 43620 34860 43920
rect 34980 43620 35010 43920
rect 35070 43620 35100 43920
rect 35940 43320 35970 43920
rect 36030 43890 36240 43920
rect 36030 43440 36060 43890
rect 36210 43440 36240 43890
rect 36030 43320 36240 43440
rect 36300 43320 36390 43920
rect 36450 43860 36750 43920
rect 36450 43440 36540 43860
rect 36660 43440 36750 43860
rect 36450 43320 36750 43440
rect 36810 43320 36900 43920
rect 36960 43890 37170 43920
rect 36960 43440 36990 43890
rect 37140 43440 37170 43890
rect 36960 43320 37170 43440
rect 37230 43320 37260 43920
rect 37860 43320 37890 43920
rect 37950 43320 37980 43920
rect 38100 43320 38130 43920
rect 38190 43890 38370 43920
rect 38190 43470 38220 43890
rect 38340 43470 38370 43890
rect 38190 43320 38370 43470
rect 38430 43320 38460 43920
rect 39540 43320 39570 43920
rect 39630 43890 39840 43920
rect 39630 43440 39660 43890
rect 39810 43440 39840 43890
rect 39630 43320 39840 43440
rect 39900 43320 39990 43920
rect 40050 43860 40350 43920
rect 40050 43440 40140 43860
rect 40260 43440 40350 43860
rect 40050 43320 40350 43440
rect 40410 43320 40500 43920
rect 40560 43890 40770 43920
rect 40560 43440 40590 43890
rect 40740 43440 40770 43890
rect 40560 43320 40770 43440
rect 40830 43320 40860 43920
rect 41940 43650 41970 43920
rect 41820 43620 41970 43650
rect 42030 43650 42060 43920
rect 42030 43620 42180 43650
rect 43140 43320 43170 43920
rect 43230 43890 43410 43920
rect 43230 43470 43260 43890
rect 43380 43470 43410 43890
rect 43230 43320 43410 43470
rect 43470 43320 43500 43920
rect 43620 43320 43650 43920
rect 43710 43320 43740 43920
rect 44340 43320 44370 43920
rect 44430 43890 44610 43920
rect 44430 43470 44460 43890
rect 44580 43470 44610 43890
rect 44430 43320 44610 43470
rect 44670 43320 44700 43920
rect 44820 43320 44850 43920
rect 44910 43320 44940 43920
rect 45300 43650 45330 43920
rect 45180 43620 45330 43650
rect 45390 43650 45420 43920
rect 45390 43620 45540 43650
rect 45780 43320 45810 43920
rect 45870 43890 46080 43920
rect 45870 43440 45900 43890
rect 46050 43440 46080 43890
rect 45870 43320 46080 43440
rect 46140 43320 46230 43920
rect 46290 43860 46590 43920
rect 46290 43440 46380 43860
rect 46500 43440 46590 43860
rect 46290 43320 46590 43440
rect 46650 43320 46740 43920
rect 46800 43890 47010 43920
rect 46800 43440 46830 43890
rect 46980 43440 47010 43890
rect 46800 43320 47010 43440
rect 47070 43320 47100 43920
rect 47460 43320 47490 43920
rect 47550 43890 47760 43920
rect 47550 43440 47580 43890
rect 47730 43440 47760 43890
rect 47550 43320 47760 43440
rect 47820 43320 47910 43920
rect 47970 43860 48270 43920
rect 47970 43440 48060 43860
rect 48180 43440 48270 43860
rect 47970 43320 48270 43440
rect 48330 43320 48420 43920
rect 48480 43890 48690 43920
rect 48480 43440 48510 43890
rect 48660 43440 48690 43890
rect 48480 43320 48690 43440
rect 48750 43320 48780 43920
rect 6030 38280 6060 38880
rect 6120 38280 6210 38880
rect 6270 38280 6300 38880
rect 6420 38280 6450 38580
rect 6510 38280 6540 38580
rect 8430 38280 8460 38880
rect 8520 38280 8610 38880
rect 8670 38280 8700 38880
rect 9780 38280 9810 38880
rect 9870 38280 9960 38880
rect 10020 38280 10050 38880
rect 10740 38280 10770 38580
rect 10830 38280 10860 38580
rect 10980 38280 11010 38880
rect 11070 38280 11160 38880
rect 11220 38280 11250 38880
rect 11700 38280 11730 38880
rect 11790 38760 12000 38880
rect 11790 38310 11820 38760
rect 11970 38310 12000 38760
rect 11790 38280 12000 38310
rect 12060 38280 12150 38880
rect 12210 38760 12510 38880
rect 12210 38340 12300 38760
rect 12420 38340 12510 38760
rect 12210 38280 12510 38340
rect 12570 38280 12660 38880
rect 12720 38760 12930 38880
rect 12720 38310 12750 38760
rect 12900 38310 12930 38760
rect 12720 38280 12930 38310
rect 12990 38280 13020 38880
rect 13620 38280 13650 38880
rect 13710 38280 13800 38880
rect 13860 38280 13890 38880
rect 14670 38280 14700 38580
rect 14760 38280 14790 38580
rect 14910 38280 14940 38880
rect 15000 38280 15090 38880
rect 15150 38280 15180 38880
rect 15660 38550 15810 38580
rect 15780 38280 15810 38550
rect 15870 38550 16020 38580
rect 15870 38280 15900 38550
rect 16500 38280 16530 38880
rect 16590 38730 16770 38880
rect 16590 38310 16620 38730
rect 16740 38310 16770 38730
rect 16590 38280 16770 38310
rect 16830 38280 16860 38880
rect 16980 38280 17010 38880
rect 17070 38280 17100 38880
rect 17700 38280 17730 38880
rect 17790 38280 17820 38880
rect 17940 38280 17970 38880
rect 18030 38730 18210 38880
rect 18030 38310 18060 38730
rect 18180 38310 18210 38730
rect 18030 38280 18210 38310
rect 18270 38280 18300 38880
rect 18540 38550 18690 38580
rect 18660 38280 18690 38550
rect 18750 38550 18900 38580
rect 18750 38280 18780 38550
rect 19380 38280 19410 38880
rect 19470 38730 19650 38880
rect 19470 38310 19500 38730
rect 19620 38310 19650 38730
rect 19470 38280 19650 38310
rect 19710 38280 19740 38880
rect 19860 38280 19890 38880
rect 19950 38280 19980 38880
rect 21150 38280 21180 38880
rect 21240 38280 21330 38880
rect 21390 38280 21420 38880
rect 22020 38280 22050 38880
rect 22110 38760 22320 38880
rect 22110 38310 22140 38760
rect 22290 38310 22320 38760
rect 22110 38280 22320 38310
rect 22380 38280 22470 38880
rect 22530 38760 22830 38880
rect 22530 38340 22620 38760
rect 22740 38340 22830 38760
rect 22530 38280 22830 38340
rect 22890 38280 22980 38880
rect 23040 38760 23250 38880
rect 23040 38310 23070 38760
rect 23220 38310 23250 38760
rect 23040 38280 23250 38310
rect 23310 38280 23340 38880
rect 23940 38280 23970 38580
rect 24030 38280 24060 38580
rect 24180 38280 24210 38580
rect 24270 38280 24300 38580
rect 24900 38280 24930 38880
rect 24990 38730 25170 38880
rect 24990 38310 25020 38730
rect 25140 38310 25170 38730
rect 24990 38280 25170 38310
rect 25230 38280 25260 38880
rect 25380 38280 25410 38880
rect 25470 38280 25500 38880
rect 26400 38280 26430 38880
rect 26490 38280 26580 38880
rect 26640 38280 26730 38880
rect 26850 38280 26940 38880
rect 27000 38280 27090 38880
rect 27150 38280 27180 38880
rect 27900 38550 28050 38580
rect 28020 38280 28050 38550
rect 28110 38550 28260 38580
rect 28110 38280 28140 38550
rect 30750 38280 30780 38880
rect 30840 38280 30930 38880
rect 30990 38280 31020 38880
rect 32190 38280 32220 38880
rect 32280 38280 32370 38880
rect 32430 38280 32460 38880
rect 33540 38280 33570 38880
rect 33630 38760 33840 38880
rect 33630 38310 33660 38760
rect 33810 38310 33840 38760
rect 33630 38280 33840 38310
rect 33900 38280 33990 38880
rect 34050 38760 34350 38880
rect 34050 38340 34140 38760
rect 34260 38340 34350 38760
rect 34050 38280 34350 38340
rect 34410 38280 34500 38880
rect 34560 38760 34770 38880
rect 34560 38310 34590 38760
rect 34740 38310 34770 38760
rect 34560 38280 34770 38310
rect 34830 38280 34860 38880
rect 36180 38280 36210 38880
rect 36270 38730 36450 38880
rect 36270 38310 36300 38730
rect 36420 38310 36450 38730
rect 36270 38280 36450 38310
rect 36510 38280 36540 38880
rect 36660 38280 36690 38880
rect 36750 38280 36780 38880
rect 37950 38280 37980 38880
rect 38040 38280 38130 38880
rect 38190 38280 38220 38880
rect 39060 38280 39090 38880
rect 39150 38730 39330 38880
rect 39150 38310 39180 38730
rect 39300 38310 39330 38730
rect 39150 38280 39330 38310
rect 39390 38280 39420 38880
rect 39540 38280 39570 38880
rect 39630 38280 39660 38880
rect 40500 38280 40530 38880
rect 40590 38280 40680 38880
rect 40740 38280 40770 38880
rect 41820 38550 41970 38580
rect 41940 38280 41970 38550
rect 42030 38550 42180 38580
rect 42030 38280 42060 38550
rect 43140 38280 43170 38880
rect 43230 38730 43410 38880
rect 43230 38310 43260 38730
rect 43380 38310 43410 38730
rect 43230 38280 43410 38310
rect 43470 38280 43500 38880
rect 43620 38280 43650 38880
rect 43710 38280 43740 38880
rect 44700 38550 44850 38580
rect 44820 38280 44850 38550
rect 44910 38550 45060 38580
rect 44910 38280 44940 38550
rect 46020 38280 46050 38880
rect 46110 38280 46140 38880
rect 46260 38280 46290 38880
rect 46350 38730 46530 38880
rect 46350 38310 46380 38730
rect 46500 38310 46530 38730
rect 46350 38280 46530 38310
rect 46590 38280 46620 38880
rect 47700 38280 47730 38880
rect 47790 38730 47970 38880
rect 47790 38310 47820 38730
rect 47940 38310 47970 38730
rect 47790 38280 47970 38310
rect 48030 38280 48060 38880
rect 48180 38280 48210 38880
rect 48270 38280 48300 38880
rect 49470 38280 49500 38880
rect 49560 38280 49650 38880
rect 49710 38280 49740 38880
rect 5790 37320 5820 37920
rect 5880 37320 5970 37920
rect 6030 37320 6060 37920
rect 7020 37890 7170 37920
rect 7140 37740 7170 37890
rect 7020 37620 7170 37740
rect 7230 37650 7260 37920
rect 7230 37620 7380 37650
rect 8340 37320 8370 37920
rect 8430 37320 8460 37920
rect 8580 37320 8610 37920
rect 8670 37890 8850 37920
rect 8670 37470 8700 37890
rect 8820 37470 8850 37890
rect 8670 37320 8850 37470
rect 8910 37320 8940 37920
rect 10980 37320 11010 37920
rect 11070 37320 11160 37920
rect 11220 37320 11250 37920
rect 12180 37320 12210 37920
rect 12270 37320 12300 37920
rect 12420 37320 12450 37920
rect 12510 37890 12690 37920
rect 12510 37470 12540 37890
rect 12660 37470 12690 37890
rect 12510 37320 12690 37470
rect 12750 37320 12780 37920
rect 15060 37320 15090 37920
rect 15150 37320 15180 37920
rect 15300 37320 15330 37920
rect 15390 37890 15570 37920
rect 15390 37470 15420 37890
rect 15540 37470 15570 37890
rect 15390 37320 15570 37470
rect 15630 37320 15660 37920
rect 16830 37620 16860 37920
rect 16920 37620 16950 37920
rect 17070 37320 17100 37920
rect 17160 37320 17250 37920
rect 17310 37320 17340 37920
rect 18180 37320 18210 37920
rect 18270 37320 18360 37920
rect 18420 37320 18450 37920
rect 19620 37320 19650 37920
rect 19710 37320 19800 37920
rect 19860 37320 19890 37920
rect 21060 37320 21090 37920
rect 21150 37320 21240 37920
rect 21300 37320 21330 37920
rect 22500 37320 22530 37920
rect 22590 37320 22680 37920
rect 22740 37320 22770 37920
rect 23940 37650 23970 37920
rect 23820 37620 23970 37650
rect 24030 37650 24060 37920
rect 24030 37620 24180 37650
rect 25230 37320 25260 37920
rect 25320 37320 25410 37920
rect 25470 37320 25500 37920
rect 26580 37320 26610 37920
rect 26670 37890 26850 37920
rect 26670 37470 26700 37890
rect 26820 37470 26850 37890
rect 26670 37320 26850 37470
rect 26910 37320 26940 37920
rect 27060 37320 27090 37920
rect 27150 37320 27180 37920
rect 28020 37320 28050 37920
rect 28110 37320 28200 37920
rect 28260 37320 28290 37920
rect 29220 37320 29250 37920
rect 29310 37320 29400 37920
rect 29460 37320 29490 37920
rect 30180 37320 30210 37920
rect 30270 37890 30450 37920
rect 30270 37470 30300 37890
rect 30420 37470 30450 37890
rect 30270 37320 30450 37470
rect 30510 37320 30540 37920
rect 30660 37320 30690 37920
rect 30750 37320 30780 37920
rect 31380 37650 31410 37920
rect 31260 37620 31410 37650
rect 31470 37650 31500 37920
rect 31470 37620 31620 37650
rect 32100 37320 32130 37920
rect 32190 37320 32220 37920
rect 32340 37320 32370 37920
rect 32430 37890 32610 37920
rect 32430 37470 32460 37890
rect 32580 37470 32610 37890
rect 32430 37320 32610 37470
rect 32670 37320 32700 37920
rect 33390 37320 33420 37920
rect 33480 37320 33570 37920
rect 33630 37320 33660 37920
rect 34740 37320 34770 37920
rect 34830 37320 34920 37920
rect 34980 37320 35010 37920
rect 35700 37320 35730 37920
rect 35790 37890 36000 37920
rect 35790 37440 35820 37890
rect 35970 37440 36000 37890
rect 35790 37320 36000 37440
rect 36060 37320 36150 37920
rect 36210 37860 36510 37920
rect 36210 37440 36300 37860
rect 36420 37440 36510 37860
rect 36210 37320 36510 37440
rect 36570 37320 36660 37920
rect 36720 37890 36930 37920
rect 36720 37440 36750 37890
rect 36900 37440 36930 37890
rect 36720 37320 36930 37440
rect 36990 37320 37020 37920
rect 39060 37650 39090 37920
rect 38940 37620 39090 37650
rect 39150 37650 39180 37920
rect 39150 37620 39300 37650
rect 40020 37320 40050 37920
rect 40110 37320 40200 37920
rect 40260 37868 40560 37920
rect 40260 37746 40350 37868
rect 40470 37746 40560 37868
rect 40260 37522 40560 37746
rect 40260 37402 40350 37522
rect 40470 37402 40560 37522
rect 40260 37320 40560 37402
rect 40620 37320 40710 37920
rect 40770 37906 40920 37920
rect 40770 37334 40800 37906
rect 41700 37650 41730 37920
rect 41580 37620 41730 37650
rect 41790 37650 41820 37920
rect 41790 37620 41940 37650
rect 42300 37906 42450 37920
rect 40770 37320 40920 37334
rect 42420 37334 42450 37906
rect 42300 37320 42450 37334
rect 42510 37906 42690 37920
rect 42510 37334 42540 37906
rect 42660 37334 42690 37906
rect 42510 37320 42690 37334
rect 42750 37890 42930 37920
rect 42750 37470 42780 37890
rect 42900 37470 42930 37890
rect 42750 37320 42930 37470
rect 42990 37906 43140 37920
rect 42990 37334 43020 37906
rect 43620 37650 43650 37920
rect 43500 37620 43650 37650
rect 43710 37650 43740 37920
rect 43710 37620 43860 37650
rect 44460 37906 44610 37920
rect 42990 37320 43140 37334
rect 44580 37334 44610 37906
rect 44460 37320 44610 37334
rect 44670 37890 44850 37920
rect 44670 37470 44700 37890
rect 44820 37470 44850 37890
rect 44670 37320 44850 37470
rect 44910 37906 45090 37920
rect 44910 37334 44940 37906
rect 45060 37334 45090 37906
rect 44910 37320 45090 37334
rect 45150 37906 45300 37920
rect 45150 37334 45180 37906
rect 45150 37320 45300 37334
rect 46140 37906 46290 37920
rect 46260 37334 46290 37906
rect 46140 37320 46290 37334
rect 46350 37320 46440 37920
rect 46500 37906 46650 37920
rect 46500 37334 46530 37906
rect 46500 37320 46650 37334
rect 47580 37906 47730 37920
rect 47700 37334 47730 37906
rect 47580 37320 47730 37334
rect 47790 37890 47970 37920
rect 47790 37470 47820 37890
rect 47940 37470 47970 37890
rect 47790 37320 47970 37470
rect 48030 37906 48210 37920
rect 48030 37334 48060 37906
rect 48180 37334 48210 37906
rect 48030 37320 48210 37334
rect 48270 37906 48420 37920
rect 48270 37334 48300 37906
rect 48270 37320 48420 37334
rect 49350 37906 49500 37920
rect 49470 37334 49500 37906
rect 49350 37320 49500 37334
rect 49560 37320 49650 37920
rect 49710 37906 49860 37920
rect 49710 37334 49740 37906
rect 49710 37320 49860 37334
rect 6540 32866 6690 32880
rect 6660 32294 6690 32866
rect 6540 32280 6690 32294
rect 6750 32866 6930 32880
rect 6750 32294 6780 32866
rect 6900 32294 6930 32866
rect 6750 32280 6930 32294
rect 6990 32730 7170 32880
rect 6990 32310 7020 32730
rect 7140 32310 7170 32730
rect 6990 32280 7170 32310
rect 7230 32866 7380 32880
rect 7230 32294 7260 32866
rect 7230 32280 7380 32294
rect 7740 32866 7890 32880
rect 7860 32294 7890 32866
rect 7740 32280 7890 32294
rect 7950 32866 8130 32880
rect 7950 32294 7980 32866
rect 8100 32294 8130 32866
rect 7950 32280 8130 32294
rect 8190 32730 8370 32880
rect 8190 32310 8220 32730
rect 8340 32310 8370 32730
rect 8190 32280 8370 32310
rect 8430 32866 8580 32880
rect 8430 32294 8460 32866
rect 8430 32280 8580 32294
rect 8940 32866 9090 32880
rect 9060 32294 9090 32866
rect 8940 32280 9090 32294
rect 9150 32746 9360 32880
rect 9150 32324 9194 32746
rect 9316 32324 9360 32746
rect 9150 32280 9360 32324
rect 9420 32280 9510 32880
rect 9570 32760 9870 32880
rect 9570 32340 9660 32760
rect 9780 32340 9870 32760
rect 9570 32280 9870 32340
rect 9930 32280 10020 32880
rect 10080 32746 10290 32880
rect 10080 32324 10124 32746
rect 10246 32324 10290 32746
rect 10080 32280 10290 32324
rect 10350 32866 10500 32880
rect 10350 32294 10380 32866
rect 10350 32280 10500 32294
rect 11100 32866 11250 32880
rect 11220 32294 11250 32866
rect 11100 32280 11250 32294
rect 11310 32746 11520 32880
rect 11310 32324 11354 32746
rect 11476 32324 11520 32746
rect 11310 32280 11520 32324
rect 11580 32280 11670 32880
rect 11730 32760 12030 32880
rect 11730 32340 11820 32760
rect 11940 32340 12030 32760
rect 11730 32280 12030 32340
rect 12090 32280 12180 32880
rect 12240 32746 12450 32880
rect 12240 32324 12284 32746
rect 12406 32324 12450 32746
rect 12240 32280 12450 32324
rect 12510 32866 12660 32880
rect 12510 32294 12540 32866
rect 15180 32866 15330 32880
rect 12510 32280 12660 32294
rect 13740 32550 13890 32580
rect 13860 32280 13890 32550
rect 13950 32550 14100 32580
rect 13950 32280 13980 32550
rect 15300 32294 15330 32866
rect 15180 32280 15330 32294
rect 15390 32280 15480 32880
rect 15540 32866 15690 32880
rect 15540 32294 15570 32866
rect 15540 32280 15690 32294
rect 16620 32866 16770 32880
rect 16740 32294 16770 32866
rect 16620 32280 16770 32294
rect 16830 32730 17010 32880
rect 16830 32310 16860 32730
rect 16980 32310 17010 32730
rect 16830 32280 17010 32310
rect 17070 32866 17250 32880
rect 17070 32294 17100 32866
rect 17220 32294 17250 32866
rect 17070 32280 17250 32294
rect 17310 32866 17460 32880
rect 17310 32294 17340 32866
rect 17310 32280 17460 32294
rect 19350 32866 19500 32880
rect 19470 32294 19500 32866
rect 19350 32280 19500 32294
rect 19560 32280 19650 32880
rect 19710 32866 19860 32880
rect 19710 32294 19740 32866
rect 21030 32866 21180 32880
rect 19710 32280 19860 32294
rect 20790 32566 20940 32580
rect 20910 32294 20940 32566
rect 20790 32280 20940 32294
rect 21000 32294 21030 32580
rect 21150 32294 21180 32866
rect 21000 32280 21180 32294
rect 21240 32280 21330 32880
rect 21390 32866 21540 32880
rect 21390 32294 21420 32866
rect 21390 32280 21540 32294
rect 23340 32866 23490 32880
rect 23460 32294 23490 32866
rect 23340 32280 23490 32294
rect 23550 32730 23730 32880
rect 23550 32310 23580 32730
rect 23700 32310 23730 32730
rect 23550 32280 23730 32310
rect 23790 32866 23970 32880
rect 23790 32294 23820 32866
rect 23940 32294 23970 32866
rect 23790 32280 23970 32294
rect 24030 32866 24180 32880
rect 24030 32294 24060 32866
rect 24030 32280 24180 32294
rect 24780 32866 24930 32880
rect 24900 32294 24930 32866
rect 24780 32280 24930 32294
rect 24990 32730 25170 32880
rect 24990 32310 25020 32730
rect 25140 32310 25170 32730
rect 24990 32280 25170 32310
rect 25230 32866 25410 32880
rect 25230 32294 25260 32866
rect 25380 32294 25410 32866
rect 25230 32280 25410 32294
rect 25470 32866 25620 32880
rect 25470 32294 25500 32866
rect 25470 32280 25620 32294
rect 25980 32866 26130 32880
rect 26100 32294 26130 32866
rect 25980 32280 26130 32294
rect 26190 32746 26400 32880
rect 26190 32324 26234 32746
rect 26356 32324 26400 32746
rect 26190 32280 26400 32324
rect 26460 32280 26550 32880
rect 26610 32760 26910 32880
rect 26610 32340 26700 32760
rect 26820 32340 26910 32760
rect 26610 32280 26910 32340
rect 26970 32280 27060 32880
rect 27120 32746 27330 32880
rect 27120 32324 27164 32746
rect 27286 32324 27330 32746
rect 27120 32280 27330 32324
rect 27390 32866 27540 32880
rect 27390 32294 27420 32866
rect 31110 32866 31260 32880
rect 27390 32280 27540 32294
rect 30300 32550 30450 32580
rect 30420 32280 30450 32550
rect 30510 32550 30660 32580
rect 30510 32280 30540 32550
rect 31230 32294 31260 32866
rect 31110 32280 31260 32294
rect 31320 32280 31410 32880
rect 31470 32866 31620 32880
rect 31470 32294 31500 32866
rect 31470 32280 31620 32294
rect 31980 32866 32130 32880
rect 32100 32294 32130 32866
rect 31980 32280 32130 32294
rect 32190 32730 32370 32880
rect 32190 32310 32220 32730
rect 32340 32310 32370 32730
rect 32190 32280 32370 32310
rect 32430 32866 32610 32880
rect 32430 32294 32460 32866
rect 32580 32294 32610 32866
rect 32430 32280 32610 32294
rect 32670 32866 32820 32880
rect 32670 32294 32700 32866
rect 32670 32280 32820 32294
rect 33180 32866 33330 32880
rect 33300 32294 33330 32866
rect 33180 32280 33330 32294
rect 33390 32280 33480 32880
rect 33540 32866 33690 32880
rect 33540 32294 33570 32866
rect 33540 32280 33690 32294
rect 34620 32866 34770 32880
rect 34740 32294 34770 32866
rect 34620 32280 34770 32294
rect 34830 32280 34920 32880
rect 34980 32866 35130 32880
rect 34980 32294 35010 32866
rect 34980 32280 35130 32294
rect 36060 32866 36210 32880
rect 36180 32294 36210 32866
rect 36060 32280 36210 32294
rect 36270 32280 36360 32880
rect 36420 32866 36570 32880
rect 36420 32294 36450 32866
rect 36420 32280 36570 32294
rect 37590 32866 37740 32880
rect 37710 32294 37740 32866
rect 37590 32280 37740 32294
rect 37800 32280 37890 32880
rect 37950 32866 38100 32880
rect 37950 32294 37980 32866
rect 37950 32280 38100 32294
rect 38940 32866 39090 32880
rect 39060 32294 39090 32866
rect 38940 32280 39090 32294
rect 39150 32280 39240 32880
rect 39300 32866 39450 32880
rect 39300 32294 39330 32866
rect 39300 32280 39450 32294
rect 40140 32866 40290 32880
rect 40260 32294 40290 32866
rect 40140 32280 40290 32294
rect 40350 32730 40530 32880
rect 40350 32310 40380 32730
rect 40500 32310 40530 32730
rect 40350 32280 40530 32310
rect 40590 32866 40770 32880
rect 40590 32294 40620 32866
rect 40740 32294 40770 32866
rect 40590 32280 40770 32294
rect 40830 32866 40980 32880
rect 40830 32294 40860 32866
rect 40830 32280 40980 32294
rect 41580 32866 41730 32880
rect 41700 32294 41730 32866
rect 41580 32280 41730 32294
rect 41790 32280 41880 32880
rect 41940 32866 42090 32880
rect 41940 32294 41970 32866
rect 41940 32280 42090 32294
rect 43020 32866 43170 32880
rect 43140 32294 43170 32866
rect 43020 32280 43170 32294
rect 43230 32730 43410 32880
rect 43230 32310 43260 32730
rect 43380 32310 43410 32730
rect 43230 32280 43410 32310
rect 43470 32866 43650 32880
rect 43470 32294 43500 32866
rect 43620 32294 43650 32866
rect 43470 32280 43650 32294
rect 43710 32866 43860 32880
rect 43710 32294 43740 32866
rect 43710 32280 43860 32294
rect 44220 32866 44370 32880
rect 44340 32294 44370 32866
rect 44220 32280 44370 32294
rect 44430 32746 44640 32880
rect 44430 32324 44474 32746
rect 44596 32324 44640 32746
rect 44430 32280 44640 32324
rect 44700 32280 44790 32880
rect 44850 32760 45150 32880
rect 44850 32340 44940 32760
rect 45060 32340 45150 32760
rect 44850 32280 45150 32340
rect 45210 32280 45300 32880
rect 45360 32746 45570 32880
rect 45360 32324 45404 32746
rect 45526 32324 45570 32746
rect 45360 32280 45570 32324
rect 45630 32866 45780 32880
rect 45630 32294 45660 32866
rect 45630 32280 45780 32294
rect 46140 32866 46290 32880
rect 46260 32294 46290 32866
rect 46140 32280 46290 32294
rect 46350 32730 46530 32880
rect 46350 32310 46380 32730
rect 46500 32310 46530 32730
rect 46350 32280 46530 32310
rect 46590 32866 46770 32880
rect 46590 32294 46620 32866
rect 46740 32294 46770 32866
rect 46590 32280 46770 32294
rect 46830 32866 46980 32880
rect 46830 32294 46860 32866
rect 46830 32280 46980 32294
rect 47670 32866 47820 32880
rect 47790 32294 47820 32866
rect 47670 32280 47820 32294
rect 47880 32280 47970 32880
rect 48030 32866 48180 32880
rect 48030 32294 48060 32866
rect 48030 32280 48180 32294
rect 49110 32866 49260 32880
rect 49230 32294 49260 32866
rect 49110 32280 49260 32294
rect 49320 32280 49410 32880
rect 49470 32866 49620 32880
rect 49470 32294 49500 32866
rect 49470 32280 49620 32294
rect 5340 31906 5490 31920
rect 5460 31334 5490 31906
rect 5340 31320 5490 31334
rect 5550 31876 5760 31920
rect 5550 31454 5594 31876
rect 5716 31454 5760 31876
rect 5550 31320 5760 31454
rect 5820 31320 5910 31920
rect 5970 31860 6270 31920
rect 5970 31440 6060 31860
rect 6180 31440 6270 31860
rect 5970 31320 6270 31440
rect 6330 31320 6420 31920
rect 6480 31876 6690 31920
rect 6480 31454 6524 31876
rect 6646 31454 6690 31876
rect 6480 31320 6690 31454
rect 6750 31906 6900 31920
rect 6750 31334 6780 31906
rect 6750 31320 6900 31334
rect 7980 31906 8130 31920
rect 8100 31334 8130 31906
rect 7980 31320 8130 31334
rect 8190 31890 8370 31920
rect 8190 31470 8220 31890
rect 8340 31470 8370 31890
rect 8190 31320 8370 31470
rect 8430 31906 8610 31920
rect 8430 31334 8460 31906
rect 8580 31334 8610 31906
rect 8430 31320 8610 31334
rect 8670 31906 8820 31920
rect 8670 31334 8700 31906
rect 8670 31320 8820 31334
rect 9750 31906 9900 31920
rect 9870 31334 9900 31906
rect 9750 31320 9900 31334
rect 9960 31320 10050 31920
rect 10110 31906 10260 31920
rect 10110 31334 10140 31906
rect 10110 31320 10260 31334
rect 11100 31906 11250 31920
rect 11220 31334 11250 31906
rect 11100 31320 11250 31334
rect 11310 31876 11520 31920
rect 11310 31454 11354 31876
rect 11476 31454 11520 31876
rect 11310 31320 11520 31454
rect 11580 31320 11670 31920
rect 11730 31860 12030 31920
rect 11730 31440 11820 31860
rect 11940 31440 12030 31860
rect 11730 31320 12030 31440
rect 12090 31320 12180 31920
rect 12240 31876 12450 31920
rect 12240 31454 12284 31876
rect 12406 31454 12450 31876
rect 12240 31320 12450 31454
rect 12510 31906 12660 31920
rect 12510 31334 12540 31906
rect 12510 31320 12660 31334
rect 14700 31906 14850 31920
rect 14820 31334 14850 31906
rect 14700 31320 14850 31334
rect 14910 31876 15120 31920
rect 14910 31454 14954 31876
rect 15076 31454 15120 31876
rect 14910 31320 15120 31454
rect 15180 31320 15270 31920
rect 15330 31860 15630 31920
rect 15330 31440 15420 31860
rect 15540 31440 15630 31860
rect 15330 31320 15630 31440
rect 15690 31320 15780 31920
rect 15840 31876 16050 31920
rect 15840 31454 15884 31876
rect 16006 31454 16050 31876
rect 15840 31320 16050 31454
rect 16110 31906 16260 31920
rect 16110 31334 16140 31906
rect 16110 31320 16260 31334
rect 17100 31906 17250 31920
rect 17220 31334 17250 31906
rect 17100 31320 17250 31334
rect 17310 31876 17520 31920
rect 17310 31454 17354 31876
rect 17476 31454 17520 31876
rect 17310 31320 17520 31454
rect 17580 31320 17670 31920
rect 17730 31860 18030 31920
rect 17730 31440 17820 31860
rect 17940 31440 18030 31860
rect 17730 31320 18030 31440
rect 18090 31320 18180 31920
rect 18240 31876 18450 31920
rect 18240 31454 18284 31876
rect 18406 31454 18450 31876
rect 18240 31320 18450 31454
rect 18510 31906 18660 31920
rect 18510 31334 18540 31906
rect 18510 31320 18660 31334
rect 19260 31906 19410 31920
rect 19380 31334 19410 31906
rect 19260 31320 19410 31334
rect 19470 31876 19680 31920
rect 19470 31454 19514 31876
rect 19636 31454 19680 31876
rect 19470 31320 19680 31454
rect 19740 31320 19830 31920
rect 19890 31860 20190 31920
rect 19890 31440 19980 31860
rect 20100 31440 20190 31860
rect 19890 31320 20190 31440
rect 20250 31320 20340 31920
rect 20400 31876 20610 31920
rect 20400 31454 20444 31876
rect 20566 31454 20610 31876
rect 20400 31320 20610 31454
rect 20670 31906 20820 31920
rect 20670 31334 20700 31906
rect 20670 31320 20820 31334
rect 21180 31906 21330 31920
rect 21300 31334 21330 31906
rect 21180 31320 21330 31334
rect 21390 31320 21480 31920
rect 21540 31906 21690 31920
rect 21540 31334 21570 31906
rect 21540 31320 21690 31334
rect 22140 31906 22290 31920
rect 22260 31334 22290 31906
rect 22140 31320 22290 31334
rect 22350 31906 22530 31920
rect 22350 31334 22380 31906
rect 22500 31334 22530 31906
rect 22350 31320 22530 31334
rect 22590 31890 22770 31920
rect 22590 31470 22620 31890
rect 22740 31470 22770 31890
rect 22590 31320 22770 31470
rect 22830 31906 22980 31920
rect 22830 31334 22860 31906
rect 23940 31650 23970 31920
rect 23820 31620 23970 31650
rect 24030 31650 24060 31920
rect 24030 31620 24180 31650
rect 24870 31906 25020 31920
rect 24990 31634 25020 31906
rect 24870 31620 25020 31634
rect 25080 31906 25260 31920
rect 25080 31620 25110 31906
rect 22830 31320 22980 31334
rect 25230 31334 25260 31906
rect 25110 31320 25260 31334
rect 25320 31320 25410 31920
rect 25470 31906 25620 31920
rect 25470 31334 25500 31906
rect 25470 31320 25620 31334
rect 25980 31906 26130 31920
rect 26100 31334 26130 31906
rect 25980 31320 26130 31334
rect 26190 31906 26370 31920
rect 26190 31334 26220 31906
rect 26340 31334 26370 31906
rect 26190 31320 26370 31334
rect 26430 31890 26610 31920
rect 26430 31470 26460 31890
rect 26580 31470 26610 31890
rect 26430 31320 26610 31470
rect 26670 31906 26820 31920
rect 26670 31334 26700 31906
rect 27300 31650 27330 31920
rect 27180 31620 27330 31650
rect 27390 31650 27420 31920
rect 27390 31620 27540 31650
rect 27750 31906 27900 31920
rect 26670 31320 26820 31334
rect 27870 31334 27900 31906
rect 27750 31320 27900 31334
rect 27960 31320 28050 31920
rect 28110 31906 28260 31920
rect 28110 31334 28140 31906
rect 28740 31650 28770 31920
rect 28620 31620 28770 31650
rect 28830 31650 28860 31920
rect 28830 31620 28980 31650
rect 29100 31906 29250 31920
rect 28110 31320 28260 31334
rect 29220 31334 29250 31906
rect 29100 31320 29250 31334
rect 29310 31906 29490 31920
rect 29310 31334 29340 31906
rect 29460 31334 29490 31906
rect 29310 31320 29490 31334
rect 29550 31890 29730 31920
rect 29550 31470 29580 31890
rect 29700 31470 29730 31890
rect 29550 31320 29730 31470
rect 29790 31906 29940 31920
rect 29790 31334 29820 31906
rect 29790 31320 29940 31334
rect 30780 31906 30930 31920
rect 30900 31334 30930 31906
rect 30780 31320 30930 31334
rect 30990 31876 31200 31920
rect 30990 31454 31034 31876
rect 31156 31454 31200 31876
rect 30990 31320 31200 31454
rect 31260 31320 31350 31920
rect 31410 31860 31710 31920
rect 31410 31440 31500 31860
rect 31620 31440 31710 31860
rect 31410 31320 31710 31440
rect 31770 31320 31860 31920
rect 31920 31876 32130 31920
rect 31920 31454 31964 31876
rect 32086 31454 32130 31876
rect 31920 31320 32130 31454
rect 32190 31906 32340 31920
rect 32190 31334 32220 31906
rect 32190 31320 32340 31334
rect 33180 31906 33330 31920
rect 33300 31334 33330 31906
rect 33180 31320 33330 31334
rect 33390 31320 33480 31920
rect 33540 31906 33690 31920
rect 33540 31334 33570 31906
rect 33540 31320 33690 31334
rect 34620 31906 34770 31920
rect 34740 31334 34770 31906
rect 34620 31320 34770 31334
rect 34830 31320 34920 31920
rect 34980 31906 35130 31920
rect 34980 31334 35010 31906
rect 34980 31320 35130 31334
rect 36060 31906 36210 31920
rect 36180 31334 36210 31906
rect 36060 31320 36210 31334
rect 36270 31906 36450 31920
rect 36270 31334 36300 31906
rect 36420 31334 36450 31906
rect 36270 31320 36450 31334
rect 36510 31890 36690 31920
rect 36510 31470 36540 31890
rect 36660 31470 36690 31890
rect 36510 31320 36690 31470
rect 36750 31906 36900 31920
rect 36750 31334 36780 31906
rect 36750 31320 36900 31334
rect 37740 31906 37890 31920
rect 37860 31334 37890 31906
rect 37740 31320 37890 31334
rect 37950 31320 38040 31920
rect 38100 31906 38250 31920
rect 38100 31334 38130 31906
rect 38100 31320 38250 31334
rect 38940 31906 39090 31920
rect 39060 31334 39090 31906
rect 38940 31320 39090 31334
rect 39150 31890 39330 31920
rect 39150 31470 39180 31890
rect 39300 31470 39330 31890
rect 39150 31320 39330 31470
rect 39390 31906 39570 31920
rect 39390 31334 39420 31906
rect 39540 31334 39570 31906
rect 39390 31320 39570 31334
rect 39630 31906 39780 31920
rect 39630 31334 39660 31906
rect 40740 31650 40770 31920
rect 40620 31620 40770 31650
rect 40830 31650 40860 31920
rect 40830 31620 40980 31650
rect 41670 31906 41820 31920
rect 39630 31320 39780 31334
rect 41790 31334 41820 31906
rect 41670 31320 41820 31334
rect 41880 31320 41970 31920
rect 42030 31906 42180 31920
rect 42030 31334 42060 31906
rect 42030 31320 42180 31334
rect 43020 31906 43170 31920
rect 43140 31334 43170 31906
rect 43020 31320 43170 31334
rect 43230 31906 43410 31920
rect 43230 31334 43260 31906
rect 43380 31334 43410 31906
rect 43230 31320 43410 31334
rect 43470 31890 43650 31920
rect 43470 31470 43500 31890
rect 43620 31470 43650 31890
rect 43470 31320 43650 31470
rect 43710 31906 43860 31920
rect 43710 31334 43740 31906
rect 43710 31320 43860 31334
rect 44460 31906 44610 31920
rect 44580 31334 44610 31906
rect 44460 31320 44610 31334
rect 44670 31890 44850 31920
rect 44670 31470 44700 31890
rect 44820 31470 44850 31890
rect 44670 31320 44850 31470
rect 44910 31906 45090 31920
rect 44910 31334 44940 31906
rect 45060 31334 45090 31906
rect 44910 31320 45090 31334
rect 45150 31906 45300 31920
rect 45150 31334 45180 31906
rect 45150 31320 45300 31334
rect 46230 31906 46380 31920
rect 46350 31334 46380 31906
rect 46230 31320 46380 31334
rect 46440 31320 46530 31920
rect 46590 31906 46740 31920
rect 46590 31334 46620 31906
rect 46590 31320 46740 31334
rect 48060 31906 48210 31920
rect 48180 31334 48210 31906
rect 48060 31320 48210 31334
rect 48270 31876 48480 31920
rect 48270 31454 48314 31876
rect 48436 31454 48480 31876
rect 48270 31320 48480 31454
rect 48540 31320 48630 31920
rect 48690 31860 48990 31920
rect 48690 31440 48780 31860
rect 48900 31440 48990 31860
rect 48690 31320 48990 31440
rect 49050 31320 49140 31920
rect 49200 31876 49410 31920
rect 49200 31454 49244 31876
rect 49366 31454 49410 31876
rect 49200 31320 49410 31454
rect 49470 31906 49620 31920
rect 49470 31334 49500 31906
rect 49470 31320 49620 31334
rect 7020 26866 7170 26880
rect 7140 26294 7170 26866
rect 7020 26280 7170 26294
rect 7230 26746 7440 26880
rect 7230 26324 7274 26746
rect 7396 26324 7440 26746
rect 7230 26280 7440 26324
rect 7500 26280 7590 26880
rect 7650 26760 7950 26880
rect 7650 26340 7740 26760
rect 7860 26340 7950 26760
rect 7650 26280 7950 26340
rect 8010 26280 8100 26880
rect 8160 26746 8370 26880
rect 8160 26324 8204 26746
rect 8326 26324 8370 26746
rect 8160 26280 8370 26324
rect 8430 26866 8580 26880
rect 8430 26294 8460 26866
rect 8430 26280 8580 26294
rect 8700 26866 8850 26880
rect 8820 26294 8850 26866
rect 8700 26280 8850 26294
rect 8910 26280 9000 26880
rect 9060 26866 9210 26880
rect 9060 26294 9090 26866
rect 9060 26280 9210 26294
rect 9420 26866 9570 26880
rect 9540 26294 9570 26866
rect 9420 26280 9570 26294
rect 9630 26746 9840 26880
rect 9630 26324 9674 26746
rect 9796 26324 9840 26746
rect 9630 26280 9840 26324
rect 9900 26280 9990 26880
rect 10050 26760 10350 26880
rect 10050 26340 10140 26760
rect 10260 26340 10350 26760
rect 10050 26280 10350 26340
rect 10410 26280 10500 26880
rect 10560 26746 10770 26880
rect 10560 26324 10604 26746
rect 10726 26324 10770 26746
rect 10560 26280 10770 26324
rect 10830 26866 10980 26880
rect 10830 26294 10860 26866
rect 10830 26280 10980 26294
rect 11100 26866 11250 26880
rect 11220 26294 11250 26866
rect 11100 26280 11250 26294
rect 11310 26730 11490 26880
rect 11310 26310 11340 26730
rect 11460 26310 11490 26730
rect 11310 26280 11490 26310
rect 11550 26866 11730 26880
rect 11550 26294 11580 26866
rect 11700 26294 11730 26866
rect 11550 26280 11730 26294
rect 11790 26866 11940 26880
rect 11790 26294 11820 26866
rect 11790 26280 11940 26294
rect 12060 26866 12210 26880
rect 12180 26294 12210 26866
rect 12060 26280 12210 26294
rect 12270 26280 12360 26880
rect 12420 26866 12570 26880
rect 12420 26294 12450 26866
rect 12420 26280 12570 26294
rect 12780 26866 12930 26880
rect 12900 26294 12930 26866
rect 12780 26280 12930 26294
rect 12990 26280 13080 26880
rect 13140 26866 13290 26880
rect 13140 26294 13170 26866
rect 14070 26866 14220 26880
rect 13140 26280 13290 26294
rect 13830 26566 13980 26580
rect 13950 26294 13980 26566
rect 13830 26280 13980 26294
rect 14040 26294 14070 26580
rect 14190 26294 14220 26866
rect 14040 26280 14220 26294
rect 14280 26280 14370 26880
rect 14430 26866 14580 26880
rect 14430 26294 14460 26866
rect 14430 26280 14580 26294
rect 15420 26866 15570 26880
rect 15540 26294 15570 26866
rect 15420 26280 15570 26294
rect 15630 26280 15720 26880
rect 15780 26866 15930 26880
rect 15780 26294 15810 26866
rect 15780 26280 15930 26294
rect 16710 26866 16860 26880
rect 16830 26294 16860 26866
rect 16710 26280 16860 26294
rect 16920 26280 17010 26880
rect 17070 26866 17220 26880
rect 17070 26294 17100 26866
rect 17070 26280 17220 26294
rect 18060 26866 18210 26880
rect 18180 26294 18210 26866
rect 18060 26280 18210 26294
rect 18270 26280 18360 26880
rect 18420 26866 18570 26880
rect 18420 26294 18450 26866
rect 18420 26280 18570 26294
rect 19260 26866 19410 26880
rect 19380 26294 19410 26866
rect 19260 26280 19410 26294
rect 19470 26866 19650 26880
rect 19470 26294 19500 26866
rect 19620 26294 19650 26866
rect 19470 26280 19650 26294
rect 19710 26730 19890 26880
rect 19710 26310 19740 26730
rect 19860 26310 19890 26730
rect 19710 26280 19890 26310
rect 19950 26866 20100 26880
rect 19950 26294 19980 26866
rect 19950 26280 20100 26294
rect 20940 26866 21090 26880
rect 21060 26294 21090 26866
rect 20940 26280 21090 26294
rect 21150 26280 21240 26880
rect 21300 26866 21450 26880
rect 21300 26294 21330 26866
rect 21300 26280 21450 26294
rect 22140 26866 22290 26880
rect 22260 26294 22290 26866
rect 22140 26280 22290 26294
rect 22350 26280 22440 26880
rect 22500 26866 22650 26880
rect 22500 26294 22530 26866
rect 22500 26280 22650 26294
rect 23580 26866 23730 26880
rect 23700 26294 23730 26866
rect 23580 26280 23730 26294
rect 23790 26280 23880 26880
rect 23940 26866 24090 26880
rect 23940 26294 23970 26866
rect 23940 26280 24090 26294
rect 25020 26866 25170 26880
rect 25140 26294 25170 26866
rect 25020 26280 25170 26294
rect 25230 26280 25320 26880
rect 25380 26866 25530 26880
rect 25380 26294 25410 26866
rect 25380 26280 25530 26294
rect 26460 26866 26610 26880
rect 26580 26294 26610 26866
rect 26460 26280 26610 26294
rect 26670 26280 26760 26880
rect 26820 26866 26970 26880
rect 26820 26294 26850 26866
rect 26820 26280 26970 26294
rect 28380 26866 28530 26880
rect 28500 26294 28530 26866
rect 28380 26280 28530 26294
rect 28590 26866 28770 26880
rect 28590 26294 28620 26866
rect 28740 26294 28770 26866
rect 28590 26280 28770 26294
rect 28830 26730 29010 26880
rect 28830 26310 28860 26730
rect 28980 26310 29010 26730
rect 28830 26280 29010 26310
rect 29070 26866 29220 26880
rect 29070 26294 29100 26866
rect 29070 26280 29220 26294
rect 30390 26866 30540 26880
rect 30510 26294 30540 26866
rect 30390 26280 30540 26294
rect 30600 26280 30690 26880
rect 30750 26866 30900 26880
rect 30750 26294 30780 26866
rect 30750 26280 30900 26294
rect 31740 26866 31890 26880
rect 31860 26294 31890 26866
rect 31740 26280 31890 26294
rect 31950 26866 32130 26880
rect 31950 26294 31980 26866
rect 32100 26294 32130 26866
rect 31950 26280 32130 26294
rect 32190 26730 32370 26880
rect 32190 26310 32220 26730
rect 32340 26310 32370 26730
rect 32190 26280 32370 26310
rect 32430 26866 32580 26880
rect 32430 26294 32460 26866
rect 32430 26280 32580 26294
rect 32940 26866 33090 26880
rect 33060 26294 33090 26866
rect 32940 26280 33090 26294
rect 33150 26746 33360 26880
rect 33150 26324 33194 26746
rect 33316 26324 33360 26746
rect 33150 26280 33360 26324
rect 33420 26280 33510 26880
rect 33570 26760 33870 26880
rect 33570 26340 33660 26760
rect 33780 26340 33870 26760
rect 33570 26280 33870 26340
rect 33930 26280 34020 26880
rect 34080 26746 34290 26880
rect 34080 26324 34124 26746
rect 34246 26324 34290 26746
rect 34080 26280 34290 26324
rect 34350 26866 34500 26880
rect 34350 26294 34380 26866
rect 34350 26280 34500 26294
rect 34860 26866 35010 26880
rect 34980 26294 35010 26866
rect 34860 26280 35010 26294
rect 35070 26280 35160 26880
rect 35220 26866 35370 26880
rect 35220 26294 35250 26866
rect 35220 26280 35370 26294
rect 36060 26866 36210 26880
rect 36180 26294 36210 26866
rect 36060 26280 36210 26294
rect 36270 26280 36360 26880
rect 36420 26866 36570 26880
rect 36420 26294 36450 26866
rect 36420 26280 36570 26294
rect 37590 26866 37740 26880
rect 37710 26294 37740 26866
rect 37590 26280 37740 26294
rect 37800 26280 37890 26880
rect 37950 26866 38100 26880
rect 37950 26294 37980 26866
rect 37950 26280 38100 26294
rect 38700 26866 38850 26880
rect 38820 26294 38850 26866
rect 38700 26280 38850 26294
rect 38910 26280 39000 26880
rect 39060 26866 39210 26880
rect 39060 26294 39090 26866
rect 39060 26280 39210 26294
rect 39660 26866 39810 26880
rect 39780 26294 39810 26866
rect 39660 26280 39810 26294
rect 39870 26746 40080 26880
rect 39870 26324 39914 26746
rect 40036 26324 40080 26746
rect 39870 26280 40080 26324
rect 40140 26280 40230 26880
rect 40290 26760 40590 26880
rect 40290 26340 40380 26760
rect 40500 26340 40590 26760
rect 40290 26280 40590 26340
rect 40650 26280 40740 26880
rect 40800 26746 41010 26880
rect 40800 26324 40844 26746
rect 40966 26324 41010 26746
rect 40800 26280 41010 26324
rect 41070 26866 41220 26880
rect 41070 26294 41100 26866
rect 41070 26280 41220 26294
rect 41580 26866 41730 26880
rect 41700 26294 41730 26866
rect 41580 26280 41730 26294
rect 41790 26280 41880 26880
rect 41940 26866 42090 26880
rect 41940 26294 41970 26866
rect 41940 26280 42090 26294
rect 43020 26866 43170 26880
rect 43140 26294 43170 26866
rect 43020 26280 43170 26294
rect 43230 26866 43410 26880
rect 43230 26294 43260 26866
rect 43380 26294 43410 26866
rect 43230 26280 43410 26294
rect 43470 26730 43650 26880
rect 43470 26310 43500 26730
rect 43620 26310 43650 26730
rect 43470 26280 43650 26310
rect 43710 26866 43860 26880
rect 43710 26294 43740 26866
rect 43710 26280 43860 26294
rect 44460 26866 44610 26880
rect 44580 26294 44610 26866
rect 44460 26280 44610 26294
rect 44670 26730 44850 26880
rect 44670 26310 44700 26730
rect 44820 26310 44850 26730
rect 44670 26280 44850 26310
rect 44910 26866 45090 26880
rect 44910 26294 44940 26866
rect 45060 26294 45090 26866
rect 44910 26280 45090 26294
rect 45150 26866 45300 26880
rect 45150 26294 45180 26866
rect 45150 26280 45300 26294
rect 45900 26866 46050 26880
rect 46020 26294 46050 26866
rect 45900 26280 46050 26294
rect 46110 26730 46290 26880
rect 46110 26310 46140 26730
rect 46260 26310 46290 26730
rect 46110 26280 46290 26310
rect 46350 26866 46530 26880
rect 46350 26294 46380 26866
rect 46500 26294 46530 26866
rect 46350 26280 46530 26294
rect 46590 26866 46740 26880
rect 46590 26294 46620 26866
rect 47340 26866 47490 26880
rect 46590 26280 46740 26294
rect 46860 26550 47010 26580
rect 46980 26280 47010 26550
rect 47070 26550 47220 26580
rect 47070 26280 47100 26550
rect 47460 26294 47490 26866
rect 47340 26280 47490 26294
rect 47550 26280 47640 26880
rect 47700 26866 48000 26880
rect 47700 26294 47790 26866
rect 47910 26294 48000 26866
rect 47700 26280 48000 26294
rect 48060 26280 48150 26880
rect 48210 26866 48360 26880
rect 48210 26294 48240 26866
rect 48210 26280 48360 26294
rect 48540 26866 48690 26880
rect 48660 26294 48690 26866
rect 48540 26280 48690 26294
rect 48750 26280 48840 26880
rect 48900 26866 49050 26880
rect 48900 26294 48930 26866
rect 48900 26280 49050 26294
rect 49260 26866 49410 26880
rect 49380 26294 49410 26866
rect 49260 26280 49410 26294
rect 49470 26730 49650 26880
rect 49470 26310 49500 26730
rect 49620 26310 49650 26730
rect 49470 26280 49650 26310
rect 49710 26866 49890 26880
rect 49710 26294 49740 26866
rect 49860 26294 49890 26866
rect 49710 26280 49890 26294
rect 49950 26866 50100 26880
rect 49950 26294 49980 26866
rect 49950 26280 50100 26294
rect 5340 25906 5490 25920
rect 5460 25334 5490 25906
rect 5340 25320 5490 25334
rect 5550 25876 5760 25920
rect 5550 25454 5594 25876
rect 5716 25454 5760 25876
rect 5550 25320 5760 25454
rect 5820 25320 5910 25920
rect 5970 25860 6270 25920
rect 5970 25440 6060 25860
rect 6180 25440 6270 25860
rect 5970 25320 6270 25440
rect 6330 25320 6420 25920
rect 6480 25876 6690 25920
rect 6480 25454 6524 25876
rect 6646 25454 6690 25876
rect 6480 25320 6690 25454
rect 6750 25906 6900 25920
rect 6750 25334 6780 25906
rect 6750 25320 6900 25334
rect 7020 25906 7170 25920
rect 7140 25334 7170 25906
rect 7020 25320 7170 25334
rect 7230 25320 7320 25920
rect 7380 25906 7530 25920
rect 7380 25334 7410 25906
rect 7380 25320 7530 25334
rect 7740 25906 7890 25920
rect 7860 25334 7890 25906
rect 7740 25320 7890 25334
rect 7950 25906 8130 25920
rect 7950 25334 7980 25906
rect 8100 25334 8130 25906
rect 7950 25320 8130 25334
rect 8190 25890 8370 25920
rect 8190 25470 8220 25890
rect 8340 25470 8370 25890
rect 8190 25320 8370 25470
rect 8430 25906 8580 25920
rect 8430 25334 8460 25906
rect 8430 25320 8580 25334
rect 8700 25906 8850 25920
rect 8820 25334 8850 25906
rect 8700 25320 8850 25334
rect 8910 25320 9000 25920
rect 9060 25906 9210 25920
rect 9060 25334 9090 25906
rect 9060 25320 9210 25334
rect 9420 25906 9570 25920
rect 9540 25334 9570 25906
rect 9420 25320 9570 25334
rect 9630 25876 9840 25920
rect 9630 25454 9674 25876
rect 9796 25454 9840 25876
rect 9630 25320 9840 25454
rect 9900 25320 9990 25920
rect 10050 25860 10350 25920
rect 10050 25440 10140 25860
rect 10260 25440 10350 25860
rect 10050 25320 10350 25440
rect 10410 25320 10500 25920
rect 10560 25876 10770 25920
rect 10560 25454 10604 25876
rect 10726 25454 10770 25876
rect 10560 25320 10770 25454
rect 10830 25906 10980 25920
rect 10830 25334 10860 25906
rect 12060 25906 12210 25920
rect 12180 25634 12210 25906
rect 12060 25620 12210 25634
rect 12270 25906 12450 25920
rect 12270 25620 12300 25906
rect 10830 25320 10980 25334
rect 12420 25334 12450 25906
rect 12300 25320 12450 25334
rect 12510 25320 12600 25920
rect 12660 25906 12810 25920
rect 12660 25334 12690 25906
rect 13860 25650 13890 25920
rect 13740 25620 13890 25650
rect 13950 25650 13980 25920
rect 13950 25620 14100 25650
rect 14940 25906 15090 25920
rect 12660 25320 12810 25334
rect 15060 25334 15090 25906
rect 14940 25320 15090 25334
rect 15150 25906 15330 25920
rect 15150 25334 15180 25906
rect 15300 25334 15330 25906
rect 15150 25320 15330 25334
rect 15390 25890 15570 25920
rect 15390 25470 15420 25890
rect 15540 25470 15570 25890
rect 15390 25320 15570 25470
rect 15630 25906 15780 25920
rect 15630 25334 15660 25906
rect 15630 25320 15780 25334
rect 20790 25906 20940 25920
rect 20910 25334 20940 25906
rect 20790 25320 20940 25334
rect 21000 25320 21090 25920
rect 21150 25906 21300 25920
rect 21150 25334 21180 25906
rect 21150 25320 21300 25334
rect 23100 25906 23250 25920
rect 23220 25334 23250 25906
rect 23100 25320 23250 25334
rect 23310 25320 23400 25920
rect 23460 25906 23610 25920
rect 23460 25334 23490 25906
rect 23460 25320 23610 25334
rect 25500 25906 25650 25920
rect 25620 25334 25650 25906
rect 25500 25320 25650 25334
rect 25710 25876 25920 25920
rect 25710 25454 25754 25876
rect 25876 25454 25920 25876
rect 25710 25320 25920 25454
rect 25980 25320 26070 25920
rect 26130 25860 26430 25920
rect 26130 25440 26220 25860
rect 26340 25440 26430 25860
rect 26130 25320 26430 25440
rect 26490 25320 26580 25920
rect 26640 25876 26850 25920
rect 26640 25454 26684 25876
rect 26806 25454 26850 25876
rect 26640 25320 26850 25454
rect 26910 25906 27060 25920
rect 26910 25334 26940 25906
rect 26910 25320 27060 25334
rect 27900 25906 28050 25920
rect 28020 25334 28050 25906
rect 27900 25320 28050 25334
rect 28110 25906 28290 25920
rect 28110 25334 28140 25906
rect 28260 25334 28290 25906
rect 28110 25320 28290 25334
rect 28350 25890 28530 25920
rect 28350 25470 28380 25890
rect 28500 25470 28530 25890
rect 28350 25320 28530 25470
rect 28590 25906 28740 25920
rect 28590 25334 28620 25906
rect 30420 25650 30450 25920
rect 30300 25620 30450 25650
rect 30510 25650 30540 25920
rect 30510 25620 30660 25650
rect 31020 25906 31170 25920
rect 28590 25320 28740 25334
rect 31140 25334 31170 25906
rect 31020 25320 31170 25334
rect 31230 25906 31410 25920
rect 31230 25334 31260 25906
rect 31380 25334 31410 25906
rect 31230 25320 31410 25334
rect 31470 25890 31650 25920
rect 31470 25470 31500 25890
rect 31620 25470 31650 25890
rect 31470 25320 31650 25470
rect 31710 25906 31860 25920
rect 31710 25334 31740 25906
rect 32340 25650 32370 25920
rect 32220 25620 32370 25650
rect 32430 25650 32460 25920
rect 32430 25620 32580 25650
rect 33180 25906 33330 25920
rect 31710 25320 31860 25334
rect 33300 25334 33330 25906
rect 33180 25320 33330 25334
rect 33390 25320 33480 25920
rect 33540 25906 33690 25920
rect 33540 25334 33570 25906
rect 33540 25320 33690 25334
rect 34620 25906 34770 25920
rect 34740 25334 34770 25906
rect 34620 25320 34770 25334
rect 34830 25320 34920 25920
rect 34980 25906 35130 25920
rect 34980 25334 35010 25906
rect 34980 25320 35130 25334
rect 36060 25906 36210 25920
rect 36180 25334 36210 25906
rect 36060 25320 36210 25334
rect 36270 25320 36360 25920
rect 36420 25906 36570 25920
rect 36420 25334 36450 25906
rect 36420 25320 36570 25334
rect 37500 25906 37650 25920
rect 37620 25334 37650 25906
rect 37500 25320 37650 25334
rect 37710 25320 37800 25920
rect 37860 25906 38010 25920
rect 37860 25334 37890 25906
rect 37860 25320 38010 25334
rect 38940 25906 39090 25920
rect 39060 25334 39090 25906
rect 38940 25320 39090 25334
rect 39150 25320 39240 25920
rect 39300 25906 39450 25920
rect 39300 25334 39330 25906
rect 39300 25320 39450 25334
rect 40380 25906 40530 25920
rect 40500 25334 40530 25906
rect 40380 25320 40530 25334
rect 40590 25320 40680 25920
rect 40740 25906 40890 25920
rect 40740 25334 40770 25906
rect 40740 25320 40890 25334
rect 41820 25906 41970 25920
rect 41940 25334 41970 25906
rect 41820 25320 41970 25334
rect 42030 25320 42120 25920
rect 42180 25906 42330 25920
rect 42180 25334 42210 25906
rect 43260 25906 43410 25920
rect 43380 25634 43410 25906
rect 43260 25620 43410 25634
rect 43470 25906 43650 25920
rect 43470 25634 43500 25906
rect 43620 25634 43650 25906
rect 43470 25620 43650 25634
rect 43710 25906 43860 25920
rect 43710 25634 43740 25906
rect 43710 25620 43860 25634
rect 44580 25650 44610 25920
rect 44460 25620 44610 25650
rect 44670 25876 44820 25920
rect 44670 25754 44700 25876
rect 44670 25620 44820 25754
rect 42180 25320 42330 25334
rect 44700 25590 44820 25620
rect 47820 25906 47970 25920
rect 47940 25334 47970 25906
rect 47820 25320 47970 25334
rect 48030 25876 48240 25920
rect 48030 25454 48074 25876
rect 48196 25454 48240 25876
rect 48030 25320 48240 25454
rect 48300 25320 48390 25920
rect 48450 25860 48750 25920
rect 48450 25440 48540 25860
rect 48660 25440 48750 25860
rect 48450 25320 48750 25440
rect 48810 25320 48900 25920
rect 48960 25876 49170 25920
rect 48960 25454 49004 25876
rect 49126 25454 49170 25876
rect 48960 25320 49170 25454
rect 49230 25906 49380 25920
rect 49230 25334 49260 25906
rect 49230 25320 49380 25334
rect 5340 20866 5490 20880
rect 5460 20294 5490 20866
rect 5340 20280 5490 20294
rect 5550 20746 5760 20880
rect 5550 20324 5594 20746
rect 5716 20324 5760 20746
rect 5550 20280 5760 20324
rect 5820 20280 5910 20880
rect 5970 20760 6270 20880
rect 5970 20340 6060 20760
rect 6180 20340 6270 20760
rect 5970 20280 6270 20340
rect 6330 20280 6420 20880
rect 6480 20746 6690 20880
rect 6480 20324 6524 20746
rect 6646 20324 6690 20746
rect 6480 20280 6690 20324
rect 6750 20866 6900 20880
rect 6750 20294 6780 20866
rect 6750 20280 6900 20294
rect 8220 20866 8370 20880
rect 8340 20294 8370 20866
rect 8220 20280 8370 20294
rect 8430 20280 8520 20880
rect 8580 20866 8730 20880
rect 8580 20294 8610 20866
rect 8580 20280 8730 20294
rect 9660 20866 9810 20880
rect 9780 20294 9810 20866
rect 9660 20280 9810 20294
rect 9870 20280 9960 20880
rect 10020 20866 10170 20880
rect 10020 20294 10050 20866
rect 10020 20280 10170 20294
rect 11100 20866 11250 20880
rect 11220 20294 11250 20866
rect 11100 20280 11250 20294
rect 11310 20866 11490 20880
rect 11310 20294 11340 20866
rect 11460 20294 11490 20866
rect 11310 20280 11490 20294
rect 11550 20730 11730 20880
rect 11550 20310 11580 20730
rect 11700 20310 11730 20730
rect 11550 20280 11730 20310
rect 11790 20866 11940 20880
rect 11790 20294 11820 20866
rect 11790 20280 11940 20294
rect 14220 20866 14370 20880
rect 14340 20294 14370 20866
rect 14220 20280 14370 20294
rect 14430 20746 14640 20880
rect 14430 20324 14474 20746
rect 14596 20324 14640 20746
rect 14430 20280 14640 20324
rect 14700 20280 14790 20880
rect 14850 20760 15150 20880
rect 14850 20340 14940 20760
rect 15060 20340 15150 20760
rect 14850 20280 15150 20340
rect 15210 20280 15300 20880
rect 15360 20746 15570 20880
rect 15360 20324 15404 20746
rect 15526 20324 15570 20746
rect 15360 20280 15570 20324
rect 15630 20866 15780 20880
rect 15630 20294 15660 20866
rect 18060 20866 18210 20880
rect 15630 20280 15780 20294
rect 16860 20446 17010 20580
rect 16980 20324 17010 20446
rect 16860 20280 17010 20324
rect 17070 20550 17220 20580
rect 17070 20280 17100 20550
rect 18180 20294 18210 20866
rect 18060 20280 18210 20294
rect 18270 20280 18360 20880
rect 18420 20866 18570 20880
rect 18420 20294 18450 20866
rect 18420 20280 18570 20294
rect 18780 20866 18930 20880
rect 18900 20294 18930 20866
rect 18780 20280 18930 20294
rect 18990 20746 19200 20880
rect 18990 20324 19034 20746
rect 19156 20324 19200 20746
rect 18990 20280 19200 20324
rect 19260 20280 19350 20880
rect 19410 20760 19710 20880
rect 19410 20340 19500 20760
rect 19620 20340 19710 20760
rect 19410 20280 19710 20340
rect 19770 20280 19860 20880
rect 19920 20746 20130 20880
rect 19920 20324 19964 20746
rect 20086 20324 20130 20746
rect 19920 20280 20130 20324
rect 20190 20866 20340 20880
rect 20190 20294 20220 20866
rect 20190 20280 20340 20294
rect 20460 20866 20610 20880
rect 20580 20294 20610 20866
rect 20460 20280 20610 20294
rect 20670 20746 20880 20880
rect 20670 20324 20714 20746
rect 20836 20324 20880 20746
rect 20670 20280 20880 20324
rect 20940 20280 21030 20880
rect 21090 20760 21390 20880
rect 21090 20340 21180 20760
rect 21300 20340 21390 20760
rect 21090 20280 21390 20340
rect 21450 20280 21540 20880
rect 21600 20746 21810 20880
rect 21600 20324 21644 20746
rect 21766 20324 21810 20746
rect 21600 20280 21810 20324
rect 21870 20866 22020 20880
rect 21870 20294 21900 20866
rect 21870 20280 22020 20294
rect 22140 20866 22290 20880
rect 22260 20294 22290 20866
rect 22140 20280 22290 20294
rect 22350 20866 22530 20880
rect 22350 20294 22380 20866
rect 22500 20294 22530 20866
rect 22350 20280 22530 20294
rect 22590 20730 22770 20880
rect 22590 20310 22620 20730
rect 22740 20310 22770 20730
rect 22590 20280 22770 20310
rect 22830 20866 22980 20880
rect 22830 20294 22860 20866
rect 26220 20866 26370 20880
rect 22830 20280 22980 20294
rect 25020 20550 25170 20580
rect 25140 20280 25170 20550
rect 25230 20550 25380 20580
rect 25230 20280 25260 20550
rect 26340 20294 26370 20866
rect 26220 20280 26370 20294
rect 26430 20866 26610 20880
rect 26430 20294 26460 20866
rect 26580 20294 26610 20866
rect 26430 20280 26610 20294
rect 26670 20730 26850 20880
rect 26670 20310 26700 20730
rect 26820 20310 26850 20730
rect 26670 20280 26850 20310
rect 26910 20866 27060 20880
rect 26910 20294 26940 20866
rect 26910 20280 27060 20294
rect 27900 20866 28050 20880
rect 28020 20294 28050 20866
rect 27900 20280 28050 20294
rect 28110 20866 28290 20880
rect 28110 20294 28140 20866
rect 28260 20294 28290 20866
rect 28110 20280 28290 20294
rect 28350 20730 28530 20880
rect 28350 20310 28380 20730
rect 28500 20310 28530 20730
rect 28350 20280 28530 20310
rect 28590 20866 28740 20880
rect 28590 20294 28620 20866
rect 28590 20280 28740 20294
rect 29100 20866 29250 20880
rect 29220 20294 29250 20866
rect 29100 20280 29250 20294
rect 29310 20280 29400 20880
rect 29460 20866 29610 20880
rect 29460 20294 29490 20866
rect 29460 20280 29610 20294
rect 30300 20866 30450 20880
rect 30420 20294 30450 20866
rect 30300 20280 30450 20294
rect 30510 20730 30690 20880
rect 30510 20310 30540 20730
rect 30660 20310 30690 20730
rect 30510 20280 30690 20310
rect 30750 20866 30930 20880
rect 30750 20294 30780 20866
rect 30900 20294 30930 20866
rect 30750 20280 30930 20294
rect 30990 20866 31140 20880
rect 30990 20294 31020 20866
rect 30990 20280 31140 20294
rect 31980 20866 32130 20880
rect 32100 20294 32130 20866
rect 31980 20280 32130 20294
rect 32190 20280 32280 20880
rect 32340 20866 32490 20880
rect 32340 20294 32370 20866
rect 32340 20280 32490 20294
rect 33180 20866 33330 20880
rect 33300 20294 33330 20866
rect 33180 20280 33330 20294
rect 33390 20280 33480 20880
rect 33540 20866 33690 20880
rect 33540 20294 33570 20866
rect 33540 20280 33690 20294
rect 34620 20866 34770 20880
rect 34740 20294 34770 20866
rect 34620 20280 34770 20294
rect 34830 20280 34920 20880
rect 34980 20866 35130 20880
rect 34980 20294 35010 20866
rect 34980 20280 35130 20294
rect 35820 20866 35970 20880
rect 35940 20294 35970 20866
rect 35820 20280 35970 20294
rect 36030 20280 36120 20880
rect 36180 20866 36330 20880
rect 36180 20294 36210 20866
rect 36180 20280 36330 20294
rect 36780 20866 36930 20880
rect 36900 20294 36930 20866
rect 36780 20280 36930 20294
rect 36990 20746 37200 20880
rect 36990 20324 37034 20746
rect 37156 20324 37200 20746
rect 36990 20280 37200 20324
rect 37260 20280 37350 20880
rect 37410 20760 37710 20880
rect 37410 20340 37500 20760
rect 37620 20340 37710 20760
rect 37410 20280 37710 20340
rect 37770 20280 37860 20880
rect 37920 20746 38130 20880
rect 37920 20324 37964 20746
rect 38086 20324 38130 20746
rect 37920 20280 38130 20324
rect 38190 20866 38340 20880
rect 38190 20294 38220 20866
rect 38190 20280 38340 20294
rect 38940 20866 39090 20880
rect 39060 20294 39090 20866
rect 38940 20280 39090 20294
rect 39150 20866 39330 20880
rect 39150 20294 39180 20866
rect 39300 20294 39330 20866
rect 39150 20280 39330 20294
rect 39390 20730 39570 20880
rect 39390 20310 39420 20730
rect 39540 20310 39570 20730
rect 39390 20280 39570 20310
rect 39630 20866 39780 20880
rect 39630 20294 39660 20866
rect 39630 20280 39780 20294
rect 40380 20866 40530 20880
rect 40500 20294 40530 20866
rect 40380 20280 40530 20294
rect 40590 20280 40680 20880
rect 40740 20866 40890 20880
rect 40740 20294 40770 20866
rect 40740 20280 40890 20294
rect 41580 20866 41730 20880
rect 41700 20294 41730 20866
rect 41580 20280 41730 20294
rect 41790 20866 41970 20880
rect 41790 20294 41820 20866
rect 41940 20294 41970 20866
rect 41790 20280 41970 20294
rect 42030 20730 42210 20880
rect 42030 20310 42060 20730
rect 42180 20310 42210 20730
rect 42030 20280 42210 20310
rect 42270 20866 42420 20880
rect 42270 20294 42300 20866
rect 44220 20866 44370 20880
rect 42270 20280 42420 20294
rect 43260 20566 43410 20580
rect 43380 20294 43410 20566
rect 43260 20280 43410 20294
rect 43470 20566 43650 20580
rect 43470 20294 43500 20566
rect 43620 20294 43650 20566
rect 43470 20280 43650 20294
rect 43710 20566 43860 20580
rect 43710 20294 43740 20566
rect 43710 20280 43860 20294
rect 44340 20294 44370 20866
rect 44220 20280 44370 20294
rect 44430 20746 44640 20880
rect 44430 20324 44474 20746
rect 44596 20324 44640 20746
rect 44430 20280 44640 20324
rect 44700 20280 44790 20880
rect 44850 20760 45150 20880
rect 44850 20340 44940 20760
rect 45060 20340 45150 20760
rect 44850 20280 45150 20340
rect 45210 20280 45300 20880
rect 45360 20746 45570 20880
rect 45360 20324 45404 20746
rect 45526 20324 45570 20746
rect 45360 20280 45570 20324
rect 45630 20866 45780 20880
rect 45630 20294 45660 20866
rect 45630 20280 45780 20294
rect 45900 20866 46050 20880
rect 46020 20294 46050 20866
rect 45900 20280 46050 20294
rect 46110 20746 46320 20880
rect 46110 20324 46154 20746
rect 46276 20324 46320 20746
rect 46110 20280 46320 20324
rect 46380 20280 46470 20880
rect 46530 20760 46830 20880
rect 46530 20340 46620 20760
rect 46740 20340 46830 20760
rect 46530 20280 46830 20340
rect 46890 20280 46980 20880
rect 47040 20746 47250 20880
rect 47040 20324 47084 20746
rect 47206 20324 47250 20746
rect 47040 20280 47250 20324
rect 47310 20866 47460 20880
rect 47310 20294 47340 20866
rect 48780 20866 48930 20880
rect 47310 20280 47460 20294
rect 47580 20550 47730 20580
rect 47700 20280 47730 20550
rect 47790 20550 47940 20580
rect 47790 20280 47820 20550
rect 48900 20294 48930 20866
rect 48780 20280 48930 20294
rect 48990 20280 49080 20880
rect 49140 20866 49440 20880
rect 49140 20294 49230 20866
rect 49350 20294 49440 20866
rect 49140 20280 49440 20294
rect 49500 20280 49590 20880
rect 49650 20866 49800 20880
rect 49650 20294 49680 20866
rect 49650 20280 49800 20294
rect 5580 19906 5730 19920
rect 5700 19334 5730 19906
rect 5580 19320 5730 19334
rect 5790 19906 5970 19920
rect 5790 19334 5820 19906
rect 5940 19334 5970 19906
rect 5790 19320 5970 19334
rect 6030 19890 6210 19920
rect 6030 19470 6060 19890
rect 6180 19470 6210 19890
rect 6030 19320 6210 19470
rect 6270 19906 6420 19920
rect 6270 19334 6300 19906
rect 6270 19320 6420 19334
rect 8940 19906 9090 19920
rect 9060 19334 9090 19906
rect 8940 19320 9090 19334
rect 9150 19876 9360 19920
rect 9150 19454 9194 19876
rect 9316 19454 9360 19876
rect 9150 19320 9360 19454
rect 9420 19320 9510 19920
rect 9570 19860 9870 19920
rect 9570 19440 9660 19860
rect 9780 19440 9870 19860
rect 9570 19320 9870 19440
rect 9930 19320 10020 19920
rect 10080 19876 10290 19920
rect 10080 19454 10124 19876
rect 10246 19454 10290 19876
rect 10080 19320 10290 19454
rect 10350 19906 10500 19920
rect 10350 19334 10380 19906
rect 10350 19320 10500 19334
rect 11580 19906 11730 19920
rect 11700 19334 11730 19906
rect 11580 19320 11730 19334
rect 11790 19876 12000 19920
rect 11790 19454 11834 19876
rect 11956 19454 12000 19876
rect 11790 19320 12000 19454
rect 12060 19320 12150 19920
rect 12210 19860 12510 19920
rect 12210 19440 12300 19860
rect 12420 19440 12510 19860
rect 12210 19320 12510 19440
rect 12570 19320 12660 19920
rect 12720 19876 12930 19920
rect 12720 19454 12764 19876
rect 12886 19454 12930 19876
rect 12720 19320 12930 19454
rect 12990 19906 13140 19920
rect 12990 19334 13020 19906
rect 12990 19320 13140 19334
rect 13500 19906 13650 19920
rect 13620 19334 13650 19906
rect 13500 19320 13650 19334
rect 13710 19876 13920 19920
rect 13710 19454 13754 19876
rect 13876 19454 13920 19876
rect 13710 19320 13920 19454
rect 13980 19320 14070 19920
rect 14130 19860 14430 19920
rect 14130 19440 14220 19860
rect 14340 19440 14430 19860
rect 14130 19320 14430 19440
rect 14490 19320 14580 19920
rect 14640 19876 14850 19920
rect 14640 19454 14684 19876
rect 14806 19454 14850 19876
rect 14640 19320 14850 19454
rect 14910 19906 15060 19920
rect 14910 19334 14940 19906
rect 14910 19320 15060 19334
rect 15510 19906 15660 19920
rect 15630 19334 15660 19906
rect 15510 19320 15660 19334
rect 15720 19320 15810 19920
rect 15870 19906 16050 19920
rect 15870 19334 15900 19906
rect 16020 19620 16050 19906
rect 16110 19906 16260 19920
rect 16110 19634 16140 19906
rect 16110 19620 16260 19634
rect 17820 19906 17970 19920
rect 15870 19320 16020 19334
rect 17940 19334 17970 19906
rect 17820 19320 17970 19334
rect 18030 19906 18210 19920
rect 18030 19334 18060 19906
rect 18180 19334 18210 19906
rect 18030 19320 18210 19334
rect 18270 19890 18450 19920
rect 18270 19470 18300 19890
rect 18420 19470 18450 19890
rect 18270 19320 18450 19470
rect 18510 19906 18660 19920
rect 18510 19334 18540 19906
rect 18510 19320 18660 19334
rect 19500 19906 19650 19920
rect 19620 19334 19650 19906
rect 19500 19320 19650 19334
rect 19710 19320 19800 19920
rect 19860 19906 20010 19920
rect 19860 19334 19890 19906
rect 19860 19320 20010 19334
rect 20940 19906 21090 19920
rect 21060 19334 21090 19906
rect 20940 19320 21090 19334
rect 21150 19320 21240 19920
rect 21300 19906 21450 19920
rect 21300 19334 21330 19906
rect 21300 19320 21450 19334
rect 22140 19906 22290 19920
rect 22260 19334 22290 19906
rect 22140 19320 22290 19334
rect 22350 19320 22440 19920
rect 22500 19906 22650 19920
rect 22500 19334 22530 19906
rect 22500 19320 22650 19334
rect 23580 19906 23730 19920
rect 23700 19334 23730 19906
rect 23580 19320 23730 19334
rect 23790 19320 23880 19920
rect 23940 19906 24090 19920
rect 23940 19334 23970 19906
rect 23940 19320 24090 19334
rect 24540 19906 24690 19920
rect 24660 19334 24690 19906
rect 24540 19320 24690 19334
rect 24750 19876 24960 19920
rect 24750 19454 24794 19876
rect 24916 19454 24960 19876
rect 24750 19320 24960 19454
rect 25020 19320 25110 19920
rect 25170 19860 25470 19920
rect 25170 19440 25260 19860
rect 25380 19440 25470 19860
rect 25170 19320 25470 19440
rect 25530 19320 25620 19920
rect 25680 19876 25890 19920
rect 25680 19454 25724 19876
rect 25846 19454 25890 19876
rect 25680 19320 25890 19454
rect 25950 19906 26100 19920
rect 25950 19334 25980 19906
rect 25950 19320 26100 19334
rect 26220 19906 26370 19920
rect 26340 19334 26370 19906
rect 26220 19320 26370 19334
rect 26430 19890 26610 19920
rect 26430 19470 26460 19890
rect 26580 19470 26610 19890
rect 26430 19320 26610 19470
rect 26670 19906 26850 19920
rect 26670 19334 26700 19906
rect 26820 19334 26850 19906
rect 26670 19320 26850 19334
rect 26910 19906 27060 19920
rect 26910 19334 26940 19906
rect 27300 19650 27330 19920
rect 27180 19620 27330 19650
rect 27390 19650 27420 19920
rect 27390 19620 27540 19650
rect 28380 19906 28530 19920
rect 26910 19320 27060 19334
rect 28500 19334 28530 19906
rect 28380 19320 28530 19334
rect 28590 19906 28770 19920
rect 28590 19334 28620 19906
rect 28740 19334 28770 19906
rect 28590 19320 28770 19334
rect 28830 19890 29010 19920
rect 28830 19470 28860 19890
rect 28980 19470 29010 19890
rect 28830 19320 29010 19470
rect 29070 19906 29220 19920
rect 29070 19334 29100 19906
rect 29070 19320 29220 19334
rect 30540 19906 30690 19920
rect 30660 19334 30690 19906
rect 30540 19320 30690 19334
rect 30750 19320 30840 19920
rect 30900 19906 31050 19920
rect 30900 19334 30930 19906
rect 30900 19320 31050 19334
rect 31980 19906 32130 19920
rect 32100 19334 32130 19906
rect 31980 19320 32130 19334
rect 32190 19320 32280 19920
rect 32340 19906 32490 19920
rect 32340 19334 32370 19906
rect 32340 19320 32490 19334
rect 33180 19906 33330 19920
rect 33300 19334 33330 19906
rect 33180 19320 33330 19334
rect 33390 19890 33570 19920
rect 33390 19470 33420 19890
rect 33540 19470 33570 19890
rect 33390 19320 33570 19470
rect 33630 19906 33810 19920
rect 33630 19334 33660 19906
rect 33780 19334 33810 19906
rect 33630 19320 33810 19334
rect 33870 19906 34020 19920
rect 33870 19334 33900 19906
rect 33870 19320 34020 19334
rect 35820 19906 35970 19920
rect 35940 19334 35970 19906
rect 35820 19320 35970 19334
rect 36030 19320 36120 19920
rect 36180 19906 36330 19920
rect 36180 19334 36210 19906
rect 36780 19906 36930 19920
rect 36900 19634 36930 19906
rect 36780 19620 36930 19634
rect 36990 19906 37170 19920
rect 36990 19620 37020 19906
rect 36180 19320 36330 19334
rect 37140 19334 37170 19906
rect 37020 19320 37170 19334
rect 37230 19320 37320 19920
rect 37380 19906 37530 19920
rect 37380 19334 37410 19906
rect 37380 19320 37530 19334
rect 37980 19906 38130 19920
rect 38100 19334 38130 19906
rect 37980 19320 38130 19334
rect 38190 19320 38280 19920
rect 38340 19906 38490 19920
rect 38340 19334 38370 19906
rect 38340 19320 38490 19334
rect 38940 19906 39090 19920
rect 39060 19334 39090 19906
rect 38940 19320 39090 19334
rect 39150 19320 39240 19920
rect 39300 19906 39450 19920
rect 39300 19334 39330 19906
rect 39300 19320 39450 19334
rect 40380 19906 40530 19920
rect 40500 19334 40530 19906
rect 40380 19320 40530 19334
rect 40590 19320 40680 19920
rect 40740 19906 40890 19920
rect 40740 19334 40770 19906
rect 41700 19650 41730 19920
rect 41580 19620 41730 19650
rect 41790 19650 41820 19920
rect 41790 19620 41940 19650
rect 42840 19906 42990 19920
rect 40740 19320 40890 19334
rect 42960 19334 42990 19906
rect 42840 19320 42990 19334
rect 43050 19320 43140 19920
rect 43200 19906 43500 19920
rect 43200 19334 43290 19906
rect 43410 19334 43500 19906
rect 43200 19320 43500 19334
rect 43560 19320 43650 19920
rect 43710 19906 43860 19920
rect 43710 19334 43740 19906
rect 43710 19320 43860 19334
rect 44460 19906 44610 19920
rect 44580 19334 44610 19906
rect 44460 19320 44610 19334
rect 44670 19890 44850 19920
rect 44670 19470 44700 19890
rect 44820 19470 44850 19890
rect 44670 19320 44850 19470
rect 44910 19906 45090 19920
rect 44910 19334 44940 19906
rect 45060 19334 45090 19906
rect 44910 19320 45090 19334
rect 45150 19906 45300 19920
rect 45150 19334 45180 19906
rect 45150 19320 45300 19334
rect 46140 19906 46290 19920
rect 46260 19334 46290 19906
rect 46140 19320 46290 19334
rect 46350 19320 46440 19920
rect 46500 19906 46650 19920
rect 46500 19334 46530 19906
rect 47580 19906 47730 19920
rect 47700 19634 47730 19906
rect 47580 19620 47730 19634
rect 47790 19906 47970 19920
rect 47790 19634 47820 19906
rect 47940 19634 47970 19906
rect 47790 19620 47970 19634
rect 48030 19906 48180 19920
rect 48030 19634 48060 19906
rect 48030 19620 48180 19634
rect 49020 19906 49170 19920
rect 46500 19320 46650 19334
rect 49140 19334 49170 19906
rect 49020 19320 49170 19334
rect 49230 19890 49410 19920
rect 49230 19470 49260 19890
rect 49380 19470 49410 19890
rect 49230 19320 49410 19470
rect 49470 19906 49650 19920
rect 49470 19334 49500 19906
rect 49620 19334 49650 19906
rect 49470 19320 49650 19334
rect 49710 19906 49860 19920
rect 49710 19334 49740 19906
rect 49710 19320 49860 19334
rect 6300 14866 6450 14880
rect 6420 14294 6450 14866
rect 6300 14280 6450 14294
rect 6510 14280 6600 14880
rect 6660 14866 6810 14880
rect 6660 14294 6690 14866
rect 6660 14280 6810 14294
rect 7740 14866 7890 14880
rect 7860 14294 7890 14866
rect 7740 14280 7890 14294
rect 7950 14746 8160 14880
rect 7950 14324 7994 14746
rect 8116 14324 8160 14746
rect 7950 14280 8160 14324
rect 8220 14280 8310 14880
rect 8370 14760 8670 14880
rect 8370 14340 8460 14760
rect 8580 14340 8670 14760
rect 8370 14280 8670 14340
rect 8730 14280 8820 14880
rect 8880 14746 9090 14880
rect 8880 14324 8924 14746
rect 9046 14324 9090 14746
rect 8880 14280 9090 14324
rect 9150 14866 9300 14880
rect 9150 14294 9180 14866
rect 9150 14280 9300 14294
rect 9420 14866 9570 14880
rect 9540 14294 9570 14866
rect 9420 14280 9570 14294
rect 9630 14746 9840 14880
rect 9630 14324 9674 14746
rect 9796 14324 9840 14746
rect 9630 14280 9840 14324
rect 9900 14280 9990 14880
rect 10050 14760 10350 14880
rect 10050 14340 10140 14760
rect 10260 14340 10350 14760
rect 10050 14280 10350 14340
rect 10410 14280 10500 14880
rect 10560 14746 10770 14880
rect 10560 14324 10604 14746
rect 10726 14324 10770 14746
rect 10560 14280 10770 14324
rect 10830 14866 10980 14880
rect 10830 14294 10860 14866
rect 10830 14280 10980 14294
rect 11100 14866 11250 14880
rect 11220 14294 11250 14866
rect 11100 14280 11250 14294
rect 11310 14746 11520 14880
rect 11310 14324 11354 14746
rect 11476 14324 11520 14746
rect 11310 14280 11520 14324
rect 11580 14280 11670 14880
rect 11730 14760 12030 14880
rect 11730 14340 11820 14760
rect 11940 14340 12030 14760
rect 11730 14280 12030 14340
rect 12090 14280 12180 14880
rect 12240 14746 12450 14880
rect 12240 14324 12284 14746
rect 12406 14324 12450 14746
rect 12240 14280 12450 14324
rect 12510 14866 12660 14880
rect 12510 14294 12540 14866
rect 12510 14280 12660 14294
rect 13260 14866 13410 14880
rect 13380 14294 13410 14866
rect 13260 14280 13410 14294
rect 13470 14746 13680 14880
rect 13470 14324 13514 14746
rect 13636 14324 13680 14746
rect 13470 14280 13680 14324
rect 13740 14280 13830 14880
rect 13890 14760 14190 14880
rect 13890 14340 13980 14760
rect 14100 14340 14190 14760
rect 13890 14280 14190 14340
rect 14250 14280 14340 14880
rect 14400 14746 14610 14880
rect 14400 14324 14444 14746
rect 14566 14324 14610 14746
rect 14400 14280 14610 14324
rect 14670 14866 14820 14880
rect 14670 14294 14700 14866
rect 14670 14280 14820 14294
rect 14940 14866 15090 14880
rect 15060 14294 15090 14866
rect 14940 14280 15090 14294
rect 15150 14746 15360 14880
rect 15150 14324 15194 14746
rect 15316 14324 15360 14746
rect 15150 14280 15360 14324
rect 15420 14280 15510 14880
rect 15570 14760 15870 14880
rect 15570 14340 15660 14760
rect 15780 14340 15870 14760
rect 15570 14280 15870 14340
rect 15930 14280 16020 14880
rect 16080 14746 16290 14880
rect 16080 14324 16124 14746
rect 16246 14324 16290 14746
rect 16080 14280 16290 14324
rect 16350 14866 16500 14880
rect 16350 14294 16380 14866
rect 16350 14280 16500 14294
rect 16710 14866 16860 14880
rect 16830 14294 16860 14866
rect 16710 14280 16860 14294
rect 16920 14280 17010 14880
rect 17070 14866 17220 14880
rect 17070 14294 17100 14866
rect 18060 14866 18210 14880
rect 17220 14294 17250 14580
rect 17070 14280 17250 14294
rect 17310 14566 17460 14580
rect 17310 14294 17340 14566
rect 17310 14280 17460 14294
rect 17580 14550 17730 14580
rect 17700 14280 17730 14550
rect 17790 14550 17940 14580
rect 17790 14280 17820 14550
rect 18180 14294 18210 14866
rect 18060 14280 18210 14294
rect 18270 14866 18450 14880
rect 18270 14294 18300 14866
rect 18420 14294 18450 14866
rect 18270 14280 18450 14294
rect 18510 14730 18690 14880
rect 18510 14310 18540 14730
rect 18660 14310 18690 14730
rect 18510 14280 18690 14310
rect 18750 14866 18900 14880
rect 18750 14294 18780 14866
rect 18750 14280 18900 14294
rect 19260 14866 19410 14880
rect 19380 14294 19410 14866
rect 19260 14280 19410 14294
rect 19470 14280 19560 14880
rect 19620 14866 19770 14880
rect 19620 14294 19650 14866
rect 19620 14280 19770 14294
rect 20700 14866 20850 14880
rect 20820 14294 20850 14866
rect 20700 14280 20850 14294
rect 20910 14730 21090 14880
rect 20910 14310 20940 14730
rect 21060 14310 21090 14730
rect 20910 14280 21090 14310
rect 21150 14866 21330 14880
rect 21150 14294 21180 14866
rect 21300 14294 21330 14866
rect 21150 14280 21330 14294
rect 21390 14866 21540 14880
rect 21390 14294 21420 14866
rect 21390 14280 21540 14294
rect 22140 14866 22290 14880
rect 22260 14294 22290 14866
rect 22140 14280 22290 14294
rect 22350 14866 22530 14880
rect 22350 14294 22380 14866
rect 22500 14294 22530 14866
rect 22350 14280 22530 14294
rect 22590 14730 22770 14880
rect 22590 14310 22620 14730
rect 22740 14310 22770 14730
rect 22590 14280 22770 14310
rect 22830 14866 22980 14880
rect 22830 14294 22860 14866
rect 22830 14280 22980 14294
rect 23580 14866 23730 14880
rect 23700 14294 23730 14866
rect 23580 14280 23730 14294
rect 23790 14280 23880 14880
rect 23940 14866 24090 14880
rect 23940 14294 23970 14866
rect 23940 14280 24090 14294
rect 24870 14866 25020 14880
rect 24990 14294 25020 14866
rect 24870 14280 25020 14294
rect 25080 14280 25170 14880
rect 25230 14866 25380 14880
rect 25230 14294 25260 14866
rect 25230 14280 25380 14294
rect 25740 14866 25890 14880
rect 25860 14294 25890 14866
rect 25740 14280 25890 14294
rect 25950 14746 26160 14880
rect 25950 14324 25994 14746
rect 26116 14324 26160 14746
rect 25950 14280 26160 14324
rect 26220 14280 26310 14880
rect 26370 14760 26670 14880
rect 26370 14340 26460 14760
rect 26580 14340 26670 14760
rect 26370 14280 26670 14340
rect 26730 14280 26820 14880
rect 26880 14746 27090 14880
rect 26880 14324 26924 14746
rect 27046 14324 27090 14746
rect 26880 14280 27090 14324
rect 27150 14866 27300 14880
rect 27150 14294 27180 14866
rect 27150 14280 27300 14294
rect 27900 14866 28050 14880
rect 28020 14294 28050 14866
rect 27900 14280 28050 14294
rect 28110 14280 28200 14880
rect 28260 14866 28410 14880
rect 28260 14294 28290 14866
rect 28260 14280 28410 14294
rect 29100 14866 29250 14880
rect 29220 14294 29250 14866
rect 29100 14280 29250 14294
rect 29310 14280 29400 14880
rect 29460 14866 29610 14880
rect 29460 14294 29490 14866
rect 29460 14280 29610 14294
rect 30300 14866 30450 14880
rect 30420 14294 30450 14866
rect 30300 14280 30450 14294
rect 30510 14746 30720 14880
rect 30510 14324 30554 14746
rect 30676 14324 30720 14746
rect 30510 14280 30720 14324
rect 30780 14280 30870 14880
rect 30930 14760 31230 14880
rect 30930 14340 31020 14760
rect 31140 14340 31230 14760
rect 30930 14280 31230 14340
rect 31290 14280 31380 14880
rect 31440 14746 31650 14880
rect 31440 14324 31484 14746
rect 31606 14324 31650 14746
rect 31440 14280 31650 14324
rect 31710 14866 31860 14880
rect 31710 14294 31740 14866
rect 31710 14280 31860 14294
rect 32310 14866 32460 14880
rect 32430 14294 32460 14866
rect 32310 14280 32460 14294
rect 32520 14280 32610 14880
rect 32670 14866 32820 14880
rect 32670 14294 32700 14866
rect 32670 14280 32820 14294
rect 33180 14866 33330 14880
rect 33300 14294 33330 14866
rect 33180 14280 33330 14294
rect 33390 14280 33480 14880
rect 33540 14866 33690 14880
rect 33540 14294 33570 14866
rect 33540 14280 33690 14294
rect 34620 14866 34770 14880
rect 34740 14294 34770 14866
rect 34620 14280 34770 14294
rect 34830 14280 34920 14880
rect 34980 14866 35130 14880
rect 34980 14294 35010 14866
rect 34980 14280 35130 14294
rect 36060 14866 36210 14880
rect 36180 14294 36210 14866
rect 36060 14280 36210 14294
rect 36270 14730 36450 14880
rect 36270 14310 36300 14730
rect 36420 14310 36450 14730
rect 36270 14280 36450 14310
rect 36510 14866 36690 14880
rect 36510 14294 36540 14866
rect 36660 14294 36690 14866
rect 36510 14280 36690 14294
rect 36750 14866 36900 14880
rect 36750 14294 36780 14866
rect 36750 14280 36900 14294
rect 37740 14866 37890 14880
rect 37860 14294 37890 14866
rect 37740 14280 37890 14294
rect 37950 14280 38040 14880
rect 38100 14866 38250 14880
rect 38100 14294 38130 14866
rect 38100 14280 38250 14294
rect 38700 14866 38850 14880
rect 38820 14294 38850 14866
rect 38700 14280 38850 14294
rect 38910 14746 39120 14880
rect 38910 14324 38954 14746
rect 39076 14324 39120 14746
rect 38910 14280 39120 14324
rect 39180 14280 39270 14880
rect 39330 14760 39630 14880
rect 39330 14340 39420 14760
rect 39540 14340 39630 14760
rect 39330 14280 39630 14340
rect 39690 14280 39780 14880
rect 39840 14746 40050 14880
rect 39840 14324 39884 14746
rect 40006 14324 40050 14746
rect 39840 14280 40050 14324
rect 40110 14866 40260 14880
rect 40110 14294 40140 14866
rect 40110 14280 40260 14294
rect 41580 14866 41730 14880
rect 41700 14294 41730 14866
rect 41580 14280 41730 14294
rect 41790 14746 42000 14880
rect 41790 14324 41834 14746
rect 41956 14324 42000 14746
rect 41790 14280 42000 14324
rect 42060 14280 42150 14880
rect 42210 14760 42510 14880
rect 42210 14340 42300 14760
rect 42420 14340 42510 14760
rect 42210 14280 42510 14340
rect 42570 14280 42660 14880
rect 42720 14746 42930 14880
rect 42720 14324 42764 14746
rect 42886 14324 42930 14746
rect 42720 14280 42930 14324
rect 42990 14866 43140 14880
rect 42990 14294 43020 14866
rect 42990 14280 43140 14294
rect 44460 14866 44610 14880
rect 44580 14294 44610 14866
rect 44460 14280 44610 14294
rect 44670 14730 44850 14880
rect 44670 14310 44700 14730
rect 44820 14310 44850 14730
rect 44670 14280 44850 14310
rect 44910 14866 45090 14880
rect 44910 14294 44940 14866
rect 45060 14294 45090 14866
rect 44910 14280 45090 14294
rect 45150 14866 45300 14880
rect 45150 14294 45180 14866
rect 45150 14280 45300 14294
rect 46140 14866 46290 14880
rect 46260 14294 46290 14866
rect 46140 14280 46290 14294
rect 46350 14280 46440 14880
rect 46500 14866 46650 14880
rect 46500 14294 46530 14866
rect 46500 14280 46650 14294
rect 47670 14866 47820 14880
rect 47790 14294 47820 14866
rect 47670 14280 47820 14294
rect 47880 14280 47970 14880
rect 48030 14866 48180 14880
rect 48030 14294 48060 14866
rect 48030 14280 48180 14294
rect 49020 14866 49170 14880
rect 49140 14294 49170 14866
rect 49020 14280 49170 14294
rect 49230 14730 49410 14880
rect 49230 14310 49260 14730
rect 49380 14310 49410 14730
rect 49230 14280 49410 14310
rect 49470 14866 49650 14880
rect 49470 14294 49500 14866
rect 49620 14294 49650 14866
rect 49470 14280 49650 14294
rect 49710 14866 49860 14880
rect 49710 14294 49740 14866
rect 49710 14280 49860 14294
rect 6870 13906 7020 13920
rect 6990 13334 7020 13906
rect 6870 13320 7020 13334
rect 7080 13320 7170 13920
rect 7230 13906 7380 13920
rect 7230 13334 7260 13906
rect 7230 13320 7380 13334
rect 8940 13906 9090 13920
rect 9060 13334 9090 13906
rect 8940 13320 9090 13334
rect 9150 13890 9330 13920
rect 9150 13470 9180 13890
rect 9300 13470 9330 13890
rect 9150 13320 9330 13470
rect 9390 13906 9570 13920
rect 9390 13334 9420 13906
rect 9540 13334 9570 13906
rect 9390 13320 9570 13334
rect 9630 13740 9810 13920
rect 9630 13320 9660 13740
rect 9780 13320 9810 13740
rect 9870 13906 10020 13920
rect 9870 13334 9900 13906
rect 9870 13320 10020 13334
rect 10860 13906 11010 13920
rect 10980 13334 11010 13906
rect 10860 13320 11010 13334
rect 11070 13320 11160 13920
rect 11220 13906 11370 13920
rect 11220 13334 11250 13906
rect 11220 13320 11370 13334
rect 12060 13906 12210 13920
rect 12180 13334 12210 13906
rect 12060 13320 12210 13334
rect 12270 13906 12450 13920
rect 12270 13334 12300 13906
rect 12420 13334 12450 13906
rect 12270 13320 12450 13334
rect 12510 13890 12690 13920
rect 12510 13470 12540 13890
rect 12660 13470 12690 13890
rect 12510 13320 12690 13470
rect 12750 13906 12900 13920
rect 12750 13334 12780 13906
rect 12750 13320 12900 13334
rect 15900 13906 16050 13920
rect 16020 13334 16050 13906
rect 15900 13320 16050 13334
rect 16110 13320 16200 13920
rect 16260 13906 16410 13920
rect 16260 13334 16290 13906
rect 16260 13320 16410 13334
rect 16620 13906 16770 13920
rect 16740 13334 16770 13906
rect 16620 13320 16770 13334
rect 16830 13906 17010 13920
rect 16830 13334 16860 13906
rect 16980 13334 17010 13906
rect 16830 13320 17010 13334
rect 17070 13890 17250 13920
rect 17070 13470 17100 13890
rect 17220 13470 17250 13890
rect 17070 13320 17250 13470
rect 17310 13906 17460 13920
rect 17310 13334 17340 13906
rect 17310 13320 17460 13334
rect 17580 13906 17730 13920
rect 17700 13334 17730 13906
rect 17580 13320 17730 13334
rect 17790 13876 18000 13920
rect 17790 13454 17834 13876
rect 17956 13454 18000 13876
rect 17790 13320 18000 13454
rect 18060 13320 18150 13920
rect 18210 13860 18510 13920
rect 18210 13440 18300 13860
rect 18420 13440 18510 13860
rect 18210 13320 18510 13440
rect 18570 13320 18660 13920
rect 18720 13876 18930 13920
rect 18720 13454 18764 13876
rect 18886 13454 18930 13876
rect 18720 13320 18930 13454
rect 18990 13906 19140 13920
rect 18990 13334 19020 13906
rect 18990 13320 19140 13334
rect 19260 13906 19410 13920
rect 19380 13334 19410 13906
rect 19260 13320 19410 13334
rect 19470 13876 19680 13920
rect 19470 13454 19514 13876
rect 19636 13454 19680 13876
rect 19470 13320 19680 13454
rect 19740 13320 19830 13920
rect 19890 13860 20190 13920
rect 19890 13440 19980 13860
rect 20100 13440 20190 13860
rect 19890 13320 20190 13440
rect 20250 13320 20340 13920
rect 20400 13876 20610 13920
rect 20400 13454 20444 13876
rect 20566 13454 20610 13876
rect 20400 13320 20610 13454
rect 20670 13906 20820 13920
rect 20670 13334 20700 13906
rect 20670 13320 20820 13334
rect 21900 13906 22050 13920
rect 22020 13334 22050 13906
rect 21900 13320 22050 13334
rect 22110 13876 22320 13920
rect 22110 13454 22154 13876
rect 22276 13454 22320 13876
rect 22110 13320 22320 13454
rect 22380 13320 22470 13920
rect 22530 13860 22830 13920
rect 22530 13440 22620 13860
rect 22740 13440 22830 13860
rect 22530 13320 22830 13440
rect 22890 13320 22980 13920
rect 23040 13876 23250 13920
rect 23040 13454 23084 13876
rect 23206 13454 23250 13876
rect 23040 13320 23250 13454
rect 23310 13906 23460 13920
rect 23310 13334 23340 13906
rect 23310 13320 23460 13334
rect 25020 13906 25170 13920
rect 25140 13334 25170 13906
rect 25020 13320 25170 13334
rect 25230 13890 25410 13920
rect 25230 13470 25260 13890
rect 25380 13470 25410 13890
rect 25230 13320 25410 13470
rect 25470 13906 25650 13920
rect 25470 13334 25500 13906
rect 25620 13334 25650 13906
rect 25470 13320 25650 13334
rect 25710 13906 25860 13920
rect 25710 13334 25740 13906
rect 25710 13320 25860 13334
rect 26700 13906 26850 13920
rect 26820 13334 26850 13906
rect 26700 13320 26850 13334
rect 26910 13320 27000 13920
rect 27060 13906 27210 13920
rect 27060 13334 27090 13906
rect 27060 13320 27210 13334
rect 29100 13906 29250 13920
rect 29220 13334 29250 13906
rect 29100 13320 29250 13334
rect 29310 13890 29490 13920
rect 29310 13470 29340 13890
rect 29460 13470 29490 13890
rect 29310 13320 29490 13470
rect 29550 13906 29730 13920
rect 29550 13334 29580 13906
rect 29700 13334 29730 13906
rect 29550 13320 29730 13334
rect 29790 13906 29940 13920
rect 29790 13334 29820 13906
rect 29790 13320 29940 13334
rect 30300 13906 30450 13920
rect 30420 13334 30450 13906
rect 30300 13320 30450 13334
rect 30510 13906 30690 13920
rect 30510 13334 30540 13906
rect 30660 13334 30690 13906
rect 30510 13320 30690 13334
rect 30750 13890 30930 13920
rect 30750 13470 30780 13890
rect 30900 13470 30930 13890
rect 30750 13320 30930 13470
rect 30990 13906 31140 13920
rect 30990 13334 31020 13906
rect 30990 13320 31140 13334
rect 32070 13906 32220 13920
rect 32190 13334 32220 13906
rect 32070 13320 32220 13334
rect 32280 13320 32370 13920
rect 32430 13906 32580 13920
rect 32430 13334 32460 13906
rect 32430 13320 32580 13334
rect 32940 13906 33090 13920
rect 33060 13334 33090 13906
rect 32940 13320 33090 13334
rect 33150 13876 33360 13920
rect 33150 13454 33194 13876
rect 33316 13454 33360 13876
rect 33150 13320 33360 13454
rect 33420 13320 33510 13920
rect 33570 13860 33870 13920
rect 33570 13440 33660 13860
rect 33780 13440 33870 13860
rect 33570 13320 33870 13440
rect 33930 13320 34020 13920
rect 34080 13876 34290 13920
rect 34080 13454 34124 13876
rect 34246 13454 34290 13876
rect 34080 13320 34290 13454
rect 34350 13906 34500 13920
rect 34350 13334 34380 13906
rect 34350 13320 34500 13334
rect 34620 13906 34770 13920
rect 34740 13334 34770 13906
rect 34620 13320 34770 13334
rect 34830 13890 35010 13920
rect 34830 13470 34860 13890
rect 34980 13470 35010 13890
rect 34830 13320 35010 13470
rect 35070 13906 35250 13920
rect 35070 13334 35100 13906
rect 35220 13334 35250 13906
rect 35070 13320 35250 13334
rect 35310 13906 35460 13920
rect 35310 13334 35340 13906
rect 35310 13320 35460 13334
rect 36060 13906 36210 13920
rect 36180 13334 36210 13906
rect 36060 13320 36210 13334
rect 36270 13320 36360 13920
rect 36420 13906 36570 13920
rect 36420 13334 36450 13906
rect 36420 13320 36570 13334
rect 37500 13906 37650 13920
rect 37620 13334 37650 13906
rect 37500 13320 37650 13334
rect 37710 13320 37800 13920
rect 37860 13906 38010 13920
rect 37860 13334 37890 13906
rect 37860 13320 38010 13334
rect 38940 13906 39090 13920
rect 39060 13334 39090 13906
rect 38940 13320 39090 13334
rect 39150 13320 39240 13920
rect 39300 13906 39450 13920
rect 39300 13334 39330 13906
rect 39300 13320 39450 13334
rect 40140 13906 40290 13920
rect 40260 13334 40290 13906
rect 40140 13320 40290 13334
rect 40350 13906 40530 13920
rect 40350 13334 40380 13906
rect 40500 13334 40530 13906
rect 40350 13320 40530 13334
rect 40590 13890 40770 13920
rect 40590 13470 40620 13890
rect 40740 13470 40770 13890
rect 40590 13320 40770 13470
rect 40830 13906 40980 13920
rect 40830 13334 40860 13906
rect 40830 13320 40980 13334
rect 41580 13906 41730 13920
rect 41700 13334 41730 13906
rect 41580 13320 41730 13334
rect 41790 13320 41880 13920
rect 41940 13906 42120 13920
rect 41940 13334 41970 13906
rect 42090 13620 42120 13906
rect 42180 13906 42330 13920
rect 42180 13634 42210 13906
rect 42180 13620 42330 13634
rect 43260 13906 43410 13920
rect 41940 13320 42090 13334
rect 43380 13334 43410 13906
rect 43260 13320 43410 13334
rect 43470 13320 43560 13920
rect 43620 13906 43770 13920
rect 43620 13334 43650 13906
rect 43620 13320 43770 13334
rect 44460 13906 44610 13920
rect 44580 13334 44610 13906
rect 44460 13320 44610 13334
rect 44670 13890 44850 13920
rect 44670 13470 44700 13890
rect 44820 13470 44850 13890
rect 44670 13320 44850 13470
rect 44910 13906 45090 13920
rect 44910 13334 44940 13906
rect 45060 13334 45090 13906
rect 44910 13320 45090 13334
rect 45150 13906 45300 13920
rect 45150 13334 45180 13906
rect 45150 13320 45300 13334
rect 46140 13906 46290 13920
rect 46260 13334 46290 13906
rect 46140 13320 46290 13334
rect 46350 13320 46440 13920
rect 46500 13906 46650 13920
rect 46500 13334 46530 13906
rect 46500 13320 46650 13334
rect 47580 13906 47730 13920
rect 47700 13334 47730 13906
rect 47580 13320 47730 13334
rect 47790 13890 47970 13920
rect 47790 13470 47820 13890
rect 47940 13470 47970 13890
rect 47790 13320 47970 13470
rect 48030 13906 48210 13920
rect 48030 13334 48060 13906
rect 48180 13334 48210 13906
rect 48030 13320 48210 13334
rect 48270 13906 48420 13920
rect 48270 13334 48300 13906
rect 48270 13320 48420 13334
rect 49350 13906 49500 13920
rect 49470 13334 49500 13906
rect 49350 13320 49500 13334
rect 49560 13320 49650 13920
rect 49710 13906 49860 13920
rect 49710 13334 49740 13906
rect 49710 13320 49860 13334
rect 5580 8866 5730 8880
rect 5700 8294 5730 8866
rect 5580 8280 5730 8294
rect 5790 8866 5970 8880
rect 5790 8294 5820 8866
rect 5940 8294 5970 8866
rect 5790 8280 5970 8294
rect 6030 8730 6210 8880
rect 6030 8310 6060 8730
rect 6180 8310 6210 8730
rect 6030 8280 6210 8310
rect 6270 8866 6420 8880
rect 6270 8294 6300 8866
rect 6270 8280 6420 8294
rect 6780 8866 6930 8880
rect 6900 8294 6930 8866
rect 6780 8280 6930 8294
rect 6990 8280 7080 8880
rect 7140 8866 7290 8880
rect 7140 8294 7170 8866
rect 7140 8280 7290 8294
rect 7740 8866 7890 8880
rect 7860 8294 7890 8866
rect 7740 8280 7890 8294
rect 7950 8746 8160 8880
rect 7950 8324 7994 8746
rect 8116 8324 8160 8746
rect 7950 8280 8160 8324
rect 8220 8280 8310 8880
rect 8370 8760 8670 8880
rect 8370 8340 8460 8760
rect 8580 8340 8670 8760
rect 8370 8280 8670 8340
rect 8730 8280 8820 8880
rect 8880 8746 9090 8880
rect 8880 8324 8924 8746
rect 9046 8324 9090 8746
rect 8880 8280 9090 8324
rect 9150 8866 9300 8880
rect 9150 8294 9180 8866
rect 9990 8866 10140 8880
rect 9150 8280 9300 8294
rect 9750 8566 9900 8580
rect 9870 8294 9900 8566
rect 9750 8280 9900 8294
rect 9960 8294 9990 8580
rect 10110 8294 10140 8866
rect 9960 8280 10140 8294
rect 10200 8280 10290 8880
rect 10350 8866 10500 8880
rect 10350 8294 10380 8866
rect 10350 8280 10500 8294
rect 11430 8866 11580 8880
rect 11550 8294 11580 8866
rect 11430 8280 11580 8294
rect 11640 8280 11730 8880
rect 11790 8866 11940 8880
rect 11790 8294 11820 8866
rect 11790 8280 11940 8294
rect 13740 8866 13890 8880
rect 13860 8294 13890 8866
rect 13740 8280 13890 8294
rect 13950 8746 14160 8880
rect 13950 8324 13994 8746
rect 14116 8324 14160 8746
rect 13950 8280 14160 8324
rect 14220 8280 14310 8880
rect 14370 8760 14670 8880
rect 14370 8340 14460 8760
rect 14580 8340 14670 8760
rect 14370 8280 14670 8340
rect 14730 8280 14820 8880
rect 14880 8746 15090 8880
rect 14880 8324 14924 8746
rect 15046 8324 15090 8746
rect 14880 8280 15090 8324
rect 15150 8866 15300 8880
rect 15150 8294 15180 8866
rect 15150 8280 15300 8294
rect 16380 8866 16530 8880
rect 16500 8294 16530 8866
rect 16380 8280 16530 8294
rect 16590 8280 16680 8880
rect 16740 8866 16890 8880
rect 16740 8294 16770 8866
rect 16740 8280 16890 8294
rect 17340 8866 17490 8880
rect 17460 8294 17490 8866
rect 17340 8280 17490 8294
rect 17550 8746 17760 8880
rect 17550 8324 17594 8746
rect 17716 8324 17760 8746
rect 17550 8280 17760 8324
rect 17820 8280 17910 8880
rect 17970 8760 18270 8880
rect 17970 8340 18060 8760
rect 18180 8340 18270 8760
rect 17970 8280 18270 8340
rect 18330 8280 18420 8880
rect 18480 8746 18690 8880
rect 18480 8324 18524 8746
rect 18646 8324 18690 8746
rect 18480 8280 18690 8324
rect 18750 8866 18900 8880
rect 18750 8294 18780 8866
rect 18750 8280 18900 8294
rect 19260 8866 19410 8880
rect 19380 8294 19410 8866
rect 19260 8280 19410 8294
rect 19470 8746 19680 8880
rect 19470 8324 19514 8746
rect 19636 8324 19680 8746
rect 19470 8280 19680 8324
rect 19740 8280 19830 8880
rect 19890 8760 20190 8880
rect 19890 8340 19980 8760
rect 20100 8340 20190 8760
rect 19890 8280 20190 8340
rect 20250 8280 20340 8880
rect 20400 8746 20610 8880
rect 20400 8324 20444 8746
rect 20566 8324 20610 8746
rect 20400 8280 20610 8324
rect 20670 8866 20820 8880
rect 20670 8294 20700 8866
rect 20670 8280 20820 8294
rect 21270 8866 21420 8880
rect 21390 8294 21420 8866
rect 21270 8280 21420 8294
rect 21480 8280 21570 8880
rect 21630 8866 21780 8880
rect 21630 8294 21660 8866
rect 21630 8280 21780 8294
rect 21900 8866 22050 8880
rect 22020 8294 22050 8866
rect 21900 8280 22050 8294
rect 22110 8746 22320 8880
rect 22110 8324 22154 8746
rect 22276 8324 22320 8746
rect 22110 8280 22320 8324
rect 22380 8280 22470 8880
rect 22530 8760 22830 8880
rect 22530 8340 22620 8760
rect 22740 8340 22830 8760
rect 22530 8280 22830 8340
rect 22890 8280 22980 8880
rect 23040 8746 23250 8880
rect 23040 8324 23084 8746
rect 23206 8324 23250 8746
rect 23040 8280 23250 8324
rect 23310 8866 23460 8880
rect 23310 8294 23340 8866
rect 23310 8280 23460 8294
rect 23820 8866 23970 8880
rect 23940 8294 23970 8866
rect 23820 8280 23970 8294
rect 24030 8280 24120 8880
rect 24180 8866 24330 8880
rect 24180 8294 24210 8866
rect 24180 8280 24330 8294
rect 25500 8866 25650 8880
rect 25620 8294 25650 8866
rect 25500 8280 25650 8294
rect 25710 8746 25920 8880
rect 25710 8324 25754 8746
rect 25876 8324 25920 8746
rect 25710 8280 25920 8324
rect 25980 8280 26070 8880
rect 26130 8760 26430 8880
rect 26130 8340 26220 8760
rect 26340 8340 26430 8760
rect 26130 8280 26430 8340
rect 26490 8280 26580 8880
rect 26640 8746 26850 8880
rect 26640 8324 26684 8746
rect 26806 8324 26850 8746
rect 26640 8280 26850 8324
rect 26910 8866 27060 8880
rect 26910 8294 26940 8866
rect 26910 8280 27060 8294
rect 27900 8866 28050 8880
rect 28020 8294 28050 8866
rect 27900 8280 28050 8294
rect 28110 8280 28200 8880
rect 28260 8866 28410 8880
rect 28260 8294 28290 8866
rect 31740 8866 31890 8880
rect 28260 8280 28410 8294
rect 29340 8550 29490 8580
rect 29460 8280 29490 8550
rect 29550 8550 29700 8580
rect 29550 8280 29580 8550
rect 30540 8550 30690 8580
rect 30660 8280 30690 8550
rect 30750 8550 30900 8580
rect 30750 8280 30780 8550
rect 31860 8294 31890 8866
rect 31740 8280 31890 8294
rect 31950 8730 32130 8880
rect 31950 8310 31980 8730
rect 32100 8310 32130 8730
rect 31950 8280 32130 8310
rect 32190 8866 32370 8880
rect 32190 8294 32220 8866
rect 32340 8294 32370 8866
rect 32190 8280 32370 8294
rect 32430 8866 32580 8880
rect 32430 8294 32460 8866
rect 32430 8280 32580 8294
rect 33180 8866 33330 8880
rect 33300 8294 33330 8866
rect 33180 8280 33330 8294
rect 33390 8746 33600 8880
rect 33390 8324 33434 8746
rect 33556 8324 33600 8746
rect 33390 8280 33600 8324
rect 33660 8280 33750 8880
rect 33810 8760 34110 8880
rect 33810 8340 33900 8760
rect 34020 8340 34110 8760
rect 33810 8280 34110 8340
rect 34170 8280 34260 8880
rect 34320 8746 34530 8880
rect 34320 8324 34364 8746
rect 34486 8324 34530 8746
rect 34320 8280 34530 8324
rect 34590 8866 34740 8880
rect 34590 8294 34620 8866
rect 35910 8866 36060 8880
rect 34590 8280 34740 8294
rect 35670 8566 35820 8580
rect 35790 8294 35820 8566
rect 35670 8280 35820 8294
rect 35880 8294 35910 8580
rect 36030 8294 36060 8866
rect 35880 8280 36060 8294
rect 36120 8280 36210 8880
rect 36270 8866 36420 8880
rect 36270 8294 36300 8866
rect 36270 8280 36420 8294
rect 36780 8866 36930 8880
rect 36900 8294 36930 8866
rect 36780 8280 36930 8294
rect 36990 8280 37080 8880
rect 37140 8866 37290 8880
rect 37140 8294 37170 8866
rect 38070 8866 38220 8880
rect 37140 8280 37290 8294
rect 37830 8566 37980 8580
rect 37950 8294 37980 8566
rect 37830 8280 37980 8294
rect 38040 8294 38070 8580
rect 38190 8294 38220 8866
rect 38040 8280 38220 8294
rect 38280 8280 38370 8880
rect 38430 8866 38580 8880
rect 38430 8294 38460 8866
rect 38430 8280 38580 8294
rect 38940 8866 39090 8880
rect 39060 8294 39090 8866
rect 38940 8280 39090 8294
rect 39150 8730 39330 8880
rect 39150 8310 39180 8730
rect 39300 8310 39330 8730
rect 39150 8280 39330 8310
rect 39390 8866 39570 8880
rect 39390 8294 39420 8866
rect 39540 8294 39570 8866
rect 39390 8280 39570 8294
rect 39630 8866 39780 8880
rect 39630 8294 39660 8866
rect 39630 8280 39780 8294
rect 40380 8866 40530 8880
rect 40500 8294 40530 8866
rect 40380 8280 40530 8294
rect 40590 8280 40680 8880
rect 40740 8866 40890 8880
rect 40740 8294 40770 8866
rect 40740 8280 40890 8294
rect 41580 8866 41730 8880
rect 41700 8294 41730 8866
rect 41580 8280 41730 8294
rect 41790 8280 41880 8880
rect 41940 8866 42090 8880
rect 41940 8294 41970 8866
rect 41940 8280 42090 8294
rect 42540 8866 42690 8880
rect 42660 8294 42690 8866
rect 42540 8280 42690 8294
rect 42750 8746 42960 8880
rect 42750 8324 42794 8746
rect 42916 8324 42960 8746
rect 42750 8280 42960 8324
rect 43020 8280 43110 8880
rect 43170 8760 43470 8880
rect 43170 8340 43260 8760
rect 43380 8340 43470 8760
rect 43170 8280 43470 8340
rect 43530 8280 43620 8880
rect 43680 8746 43890 8880
rect 43680 8324 43724 8746
rect 43846 8324 43890 8746
rect 43680 8280 43890 8324
rect 43950 8866 44100 8880
rect 43950 8294 43980 8866
rect 43950 8280 44100 8294
rect 45180 8866 45330 8880
rect 45300 8294 45330 8866
rect 45180 8280 45330 8294
rect 45390 8746 45600 8880
rect 45390 8324 45434 8746
rect 45556 8324 45600 8746
rect 45390 8280 45600 8324
rect 45660 8280 45750 8880
rect 45810 8760 46110 8880
rect 45810 8340 45900 8760
rect 46020 8340 46110 8760
rect 45810 8280 46110 8340
rect 46170 8280 46260 8880
rect 46320 8746 46530 8880
rect 46320 8324 46364 8746
rect 46486 8324 46530 8746
rect 46320 8280 46530 8324
rect 46590 8866 46740 8880
rect 46590 8294 46620 8866
rect 46590 8280 46740 8294
rect 47670 8866 47820 8880
rect 47790 8294 47820 8866
rect 47670 8280 47820 8294
rect 47880 8280 47970 8880
rect 48030 8866 48180 8880
rect 48030 8294 48060 8866
rect 48030 8280 48180 8294
rect 49110 8866 49260 8880
rect 49230 8294 49260 8866
rect 49110 8280 49260 8294
rect 49320 8280 49410 8880
rect 49470 8866 49620 8880
rect 49470 8294 49500 8866
rect 49470 8280 49620 8294
rect 5580 7906 5730 7920
rect 5700 7334 5730 7906
rect 5580 7320 5730 7334
rect 5790 7876 6000 7920
rect 5790 7454 5834 7876
rect 5956 7454 6000 7876
rect 5790 7320 6000 7454
rect 6060 7320 6150 7920
rect 6210 7860 6510 7920
rect 6210 7440 6300 7860
rect 6420 7440 6510 7860
rect 6210 7320 6510 7440
rect 6570 7320 6660 7920
rect 6720 7876 6930 7920
rect 6720 7454 6764 7876
rect 6886 7454 6930 7876
rect 6720 7320 6930 7454
rect 6990 7906 7140 7920
rect 6990 7334 7020 7906
rect 8100 7650 8130 7920
rect 7980 7620 8130 7650
rect 8190 7650 8220 7920
rect 8190 7620 8340 7650
rect 8700 7906 8850 7920
rect 6990 7320 7140 7334
rect 8820 7334 8850 7906
rect 8700 7320 8850 7334
rect 8910 7906 9090 7920
rect 8910 7334 8940 7906
rect 9060 7334 9090 7906
rect 8910 7320 9090 7334
rect 9150 7890 9330 7920
rect 9150 7470 9180 7890
rect 9300 7470 9330 7890
rect 9150 7320 9330 7470
rect 9390 7906 9540 7920
rect 9390 7334 9420 7906
rect 9390 7320 9540 7334
rect 9900 7906 10050 7920
rect 10020 7334 10050 7906
rect 9900 7320 10050 7334
rect 10110 7320 10200 7920
rect 10260 7906 10410 7920
rect 10260 7334 10290 7906
rect 10260 7320 10410 7334
rect 10860 7906 11010 7920
rect 10980 7334 11010 7906
rect 10860 7320 11010 7334
rect 11070 7906 11250 7920
rect 11070 7334 11100 7906
rect 11220 7334 11250 7906
rect 11070 7320 11250 7334
rect 11310 7890 11490 7920
rect 11310 7470 11340 7890
rect 11460 7470 11490 7890
rect 11310 7320 11490 7470
rect 11550 7906 11700 7920
rect 11550 7334 11580 7906
rect 11550 7320 11700 7334
rect 12300 7906 12450 7920
rect 12420 7334 12450 7906
rect 12300 7320 12450 7334
rect 12510 7320 12600 7920
rect 12660 7906 12810 7920
rect 12660 7334 12690 7906
rect 12660 7320 12810 7334
rect 13830 7906 13980 7920
rect 13950 7334 13980 7906
rect 13830 7320 13980 7334
rect 14040 7320 14130 7920
rect 14190 7906 14370 7920
rect 14190 7334 14220 7906
rect 14340 7620 14370 7906
rect 14430 7906 14580 7920
rect 14430 7634 14460 7906
rect 14430 7620 14580 7634
rect 15420 7906 15570 7920
rect 15540 7634 15570 7906
rect 15420 7620 15570 7634
rect 15630 7906 15810 7920
rect 15630 7634 15660 7906
rect 15780 7634 15810 7906
rect 15630 7620 15810 7634
rect 15870 7906 16020 7920
rect 15870 7634 15900 7906
rect 15870 7620 16020 7634
rect 18060 7906 18210 7920
rect 18180 7634 18210 7906
rect 18060 7620 18210 7634
rect 18270 7906 18450 7920
rect 18270 7634 18300 7906
rect 18420 7634 18450 7906
rect 18270 7620 18450 7634
rect 18510 7906 18660 7920
rect 18510 7634 18540 7906
rect 18510 7620 18660 7634
rect 20700 7906 20850 7920
rect 14190 7320 14340 7334
rect 20820 7334 20850 7906
rect 20700 7320 20850 7334
rect 20910 7320 21000 7920
rect 21060 7906 21210 7920
rect 21060 7334 21090 7906
rect 21060 7320 21210 7334
rect 23340 7906 23490 7920
rect 23460 7334 23490 7906
rect 23340 7320 23490 7334
rect 23550 7320 23640 7920
rect 23700 7906 23850 7920
rect 23700 7334 23730 7906
rect 23700 7320 23850 7334
rect 25740 7906 25890 7920
rect 25860 7334 25890 7906
rect 25740 7320 25890 7334
rect 25950 7876 26160 7920
rect 25950 7454 25994 7876
rect 26116 7454 26160 7876
rect 25950 7320 26160 7454
rect 26220 7320 26310 7920
rect 26370 7860 26670 7920
rect 26370 7440 26460 7860
rect 26580 7440 26670 7860
rect 26370 7320 26670 7440
rect 26730 7320 26820 7920
rect 26880 7876 27090 7920
rect 26880 7454 26924 7876
rect 27046 7454 27090 7876
rect 26880 7320 27090 7454
rect 27150 7906 27300 7920
rect 27150 7334 27180 7906
rect 27150 7320 27300 7334
rect 27900 7906 28050 7920
rect 28020 7334 28050 7906
rect 27900 7320 28050 7334
rect 28110 7320 28200 7920
rect 28260 7906 28410 7920
rect 28260 7334 28290 7906
rect 28260 7320 28410 7334
rect 29100 7906 29250 7920
rect 29220 7334 29250 7906
rect 29100 7320 29250 7334
rect 29310 7320 29400 7920
rect 29460 7906 29610 7920
rect 29460 7334 29490 7906
rect 29460 7320 29610 7334
rect 30060 7906 30210 7920
rect 30180 7334 30210 7906
rect 30060 7320 30210 7334
rect 30270 7876 30480 7920
rect 30270 7454 30314 7876
rect 30436 7454 30480 7876
rect 30270 7320 30480 7454
rect 30540 7320 30630 7920
rect 30690 7860 30990 7920
rect 30690 7440 30780 7860
rect 30900 7440 30990 7860
rect 30690 7320 30990 7440
rect 31050 7320 31140 7920
rect 31200 7876 31410 7920
rect 31200 7454 31244 7876
rect 31366 7454 31410 7876
rect 31200 7320 31410 7454
rect 31470 7906 31620 7920
rect 31470 7334 31500 7906
rect 31470 7320 31620 7334
rect 31980 7906 32130 7920
rect 32100 7334 32130 7906
rect 31980 7320 32130 7334
rect 32190 7890 32370 7920
rect 32190 7470 32220 7890
rect 32340 7470 32370 7890
rect 32190 7320 32370 7470
rect 32430 7906 32610 7920
rect 32430 7334 32460 7906
rect 32580 7334 32610 7906
rect 32430 7320 32610 7334
rect 32670 7906 32820 7920
rect 32670 7334 32700 7906
rect 32670 7320 32820 7334
rect 33180 7906 33330 7920
rect 33300 7334 33330 7906
rect 33180 7320 33330 7334
rect 33390 7320 33480 7920
rect 33540 7906 33690 7920
rect 33540 7334 33570 7906
rect 33540 7320 33690 7334
rect 34710 7906 34860 7920
rect 34830 7334 34860 7906
rect 34710 7320 34860 7334
rect 34920 7320 35010 7920
rect 35070 7906 35220 7920
rect 35070 7334 35100 7906
rect 35070 7320 35220 7334
rect 36060 7906 36210 7920
rect 36180 7334 36210 7906
rect 36060 7320 36210 7334
rect 36270 7320 36360 7920
rect 36420 7906 36570 7920
rect 36420 7334 36450 7906
rect 36420 7320 36570 7334
rect 37500 7906 37650 7920
rect 37620 7334 37650 7906
rect 37500 7320 37650 7334
rect 37710 7906 37890 7920
rect 37710 7334 37740 7906
rect 37860 7334 37890 7906
rect 37710 7320 37890 7334
rect 37950 7890 38130 7920
rect 37950 7470 37980 7890
rect 38100 7470 38130 7890
rect 37950 7320 38130 7470
rect 38190 7906 38340 7920
rect 38190 7334 38220 7906
rect 38190 7320 38340 7334
rect 38940 7906 39090 7920
rect 39060 7334 39090 7906
rect 38940 7320 39090 7334
rect 39150 7320 39240 7920
rect 39300 7906 39450 7920
rect 39300 7334 39330 7906
rect 39300 7320 39450 7334
rect 40380 7906 40530 7920
rect 40500 7334 40530 7906
rect 40380 7320 40530 7334
rect 40590 7320 40680 7920
rect 40740 7906 40890 7920
rect 40740 7334 40770 7906
rect 43260 7906 43410 7920
rect 43380 7634 43410 7906
rect 43260 7620 43410 7634
rect 43470 7906 43650 7920
rect 43470 7634 43500 7906
rect 43620 7634 43650 7906
rect 43470 7620 43650 7634
rect 43710 7906 43860 7920
rect 43710 7634 43740 7906
rect 43710 7620 43860 7634
rect 44520 7906 44670 7920
rect 40740 7320 40890 7334
rect 44640 7334 44670 7906
rect 44520 7320 44670 7334
rect 44730 7320 44820 7920
rect 44880 7906 45180 7920
rect 44880 7334 44970 7906
rect 45090 7334 45180 7906
rect 44880 7320 45180 7334
rect 45240 7320 45330 7920
rect 45390 7906 45540 7920
rect 45390 7334 45420 7906
rect 46500 7650 46530 7920
rect 46380 7620 46530 7650
rect 46590 7650 46620 7920
rect 46590 7620 46740 7650
rect 47340 7906 47490 7920
rect 45390 7320 45540 7334
rect 47460 7334 47490 7906
rect 47340 7320 47490 7334
rect 47550 7906 47730 7920
rect 47550 7334 47580 7906
rect 47700 7334 47730 7906
rect 47550 7320 47730 7334
rect 47790 7890 47970 7920
rect 47790 7470 47820 7890
rect 47940 7470 47970 7890
rect 47790 7320 47970 7470
rect 48030 7906 48180 7920
rect 48030 7334 48060 7906
rect 48030 7320 48180 7334
<< pdiffusion >>
rect 5910 42466 6060 42480
rect 5670 41866 5820 41880
rect 5790 41294 5820 41866
rect 5670 41280 5820 41294
rect 5880 41294 5910 41880
rect 6030 41294 6060 42466
rect 5880 41280 6060 41294
rect 6120 41280 6210 42480
rect 6270 42466 6420 42480
rect 6270 41294 6300 42466
rect 8070 42466 8220 42480
rect 6270 41280 6420 41294
rect 6780 41866 6930 41880
rect 6900 41294 6930 41866
rect 6780 41280 6930 41294
rect 6990 41866 7170 41880
rect 6990 41294 7020 41866
rect 7140 41294 7170 41866
rect 6990 41280 7170 41294
rect 7230 41866 7380 41880
rect 7230 41294 7260 41866
rect 7230 41280 7380 41294
rect 7830 41866 7980 41880
rect 7950 41294 7980 41866
rect 7830 41280 7980 41294
rect 8040 41294 8070 41880
rect 8190 41294 8220 42466
rect 8040 41280 8220 41294
rect 8280 41280 8370 42480
rect 8430 42466 8580 42480
rect 8430 41294 8460 42466
rect 8430 41280 8580 41294
rect 8940 42466 9090 42480
rect 9060 41294 9090 42466
rect 8940 41280 9090 41294
rect 9150 42210 9360 42480
rect 9150 41340 9194 42210
rect 9316 41340 9360 42210
rect 9150 41280 9360 41340
rect 9420 41280 9510 42480
rect 9570 42466 9870 42480
rect 9570 41294 9660 42466
rect 9780 41294 9870 42466
rect 9570 41280 9870 41294
rect 9930 41280 10020 42480
rect 10080 42210 10290 42480
rect 10080 41340 10124 42210
rect 10246 41340 10290 42210
rect 10080 41280 10290 41340
rect 10350 42466 10500 42480
rect 10350 41294 10380 42466
rect 10350 41280 10500 41294
rect 11070 41310 11100 42480
rect 10950 41280 11100 41310
rect 11160 41280 11250 42480
rect 11310 41310 11340 42480
rect 11310 41280 11460 41310
rect 12510 41310 12540 42480
rect 12390 41280 12540 41310
rect 12600 41280 12690 42480
rect 12750 41310 12780 42480
rect 12750 41280 12900 41310
rect 13740 42466 13890 42480
rect 13860 41294 13890 42466
rect 13740 41280 13890 41294
rect 13950 41280 14040 42480
rect 14100 42466 14250 42480
rect 14100 41294 14130 42466
rect 17100 42466 17250 42480
rect 14250 41294 14280 41880
rect 14100 41280 14280 41294
rect 14340 41866 14490 41880
rect 14340 41294 14370 41866
rect 14340 41280 14490 41294
rect 15420 41866 15570 41880
rect 15540 41294 15570 41866
rect 15420 41280 15570 41294
rect 15630 41866 15810 41880
rect 15630 41294 15660 41866
rect 15780 41294 15810 41866
rect 15630 41280 15810 41294
rect 15870 41866 16020 41880
rect 15870 41294 15900 41866
rect 15870 41280 16020 41294
rect 17220 41294 17250 42466
rect 17100 41280 17250 41294
rect 17310 41280 17400 42480
rect 17460 42466 17610 42480
rect 17460 41294 17490 42466
rect 19260 42466 19410 42480
rect 17610 41294 17640 41880
rect 17460 41280 17640 41294
rect 17700 41866 17850 41880
rect 17700 41294 17730 41866
rect 17700 41280 17850 41294
rect 19380 41294 19410 42466
rect 19260 41280 19410 41294
rect 19470 42210 19680 42480
rect 19470 41340 19514 42210
rect 19636 41340 19680 42210
rect 19470 41280 19680 41340
rect 19740 41280 19830 42480
rect 19890 42466 20190 42480
rect 19890 41294 19980 42466
rect 20100 41294 20190 42466
rect 19890 41280 20190 41294
rect 20250 41280 20340 42480
rect 20400 42210 20610 42480
rect 20400 41340 20444 42210
rect 20566 41340 20610 42210
rect 20400 41280 20610 41340
rect 20670 42466 20820 42480
rect 20670 41294 20700 42466
rect 22620 42466 22770 42480
rect 20670 41280 20820 41294
rect 21300 41310 21330 41880
rect 21180 41280 21330 41310
rect 21390 41310 21420 41880
rect 21390 41280 21540 41310
rect 22740 41294 22770 42466
rect 22620 41280 22770 41294
rect 22830 42210 23040 42480
rect 22830 41340 22874 42210
rect 22996 41340 23040 42210
rect 22830 41280 23040 41340
rect 23100 41280 23190 42480
rect 23250 42466 23550 42480
rect 23250 41294 23340 42466
rect 23460 41294 23550 42466
rect 23250 41280 23550 41294
rect 23610 41280 23700 42480
rect 23760 42210 23970 42480
rect 23760 41340 23804 42210
rect 23926 41340 23970 42210
rect 23760 41280 23970 41340
rect 24030 42466 24180 42480
rect 24030 41294 24060 42466
rect 25350 42466 25500 42480
rect 24030 41280 24180 41294
rect 25110 41866 25260 41880
rect 25230 41294 25260 41866
rect 25110 41280 25260 41294
rect 25320 41294 25350 41880
rect 25470 41294 25500 42466
rect 25320 41280 25500 41294
rect 25560 41280 25650 42480
rect 25710 42466 25860 42480
rect 25710 41294 25740 42466
rect 27900 42466 28050 42480
rect 25710 41280 25860 41294
rect 26700 41866 26850 41880
rect 26820 41294 26850 41866
rect 26700 41280 26850 41294
rect 26910 41866 27090 41880
rect 26910 41294 26940 41866
rect 27060 41294 27090 41866
rect 26910 41280 27090 41294
rect 27150 41866 27300 41880
rect 27150 41294 27180 41866
rect 27150 41280 27300 41294
rect 28020 41294 28050 42466
rect 27900 41280 28050 41294
rect 28110 41280 28200 42480
rect 28260 42466 28410 42480
rect 28260 41294 28290 42466
rect 30300 42466 30450 42480
rect 28410 41294 28440 41880
rect 28260 41280 28440 41294
rect 28500 41866 28650 41880
rect 28500 41294 28530 41866
rect 28500 41280 28650 41294
rect 29100 41866 29250 41880
rect 29220 41294 29250 41866
rect 29100 41280 29250 41294
rect 29310 41866 29490 41880
rect 29310 41294 29340 41866
rect 29460 41294 29490 41866
rect 29310 41280 29490 41294
rect 29550 41866 29700 41880
rect 29550 41294 29580 41866
rect 29550 41280 29700 41294
rect 30420 41294 30450 42466
rect 30300 41280 30450 41294
rect 30510 41280 30600 42480
rect 30660 42466 30810 42480
rect 30660 41294 30690 42466
rect 31740 42466 31890 42480
rect 30810 41294 30840 41880
rect 30660 41280 30840 41294
rect 30900 41866 31050 41880
rect 30900 41294 30930 41866
rect 30900 41280 31050 41294
rect 31860 41294 31890 42466
rect 31740 41280 31890 41294
rect 31950 41280 32040 42480
rect 32100 42466 32250 42480
rect 32100 41294 32130 42466
rect 32250 41294 32280 41880
rect 32100 41280 32280 41294
rect 32340 41866 32490 41880
rect 32340 41294 32370 41866
rect 32340 41280 32490 41294
rect 33180 41866 33330 41880
rect 33300 41294 33330 41866
rect 33180 41280 33330 41294
rect 33390 41866 33570 41880
rect 33390 41294 33420 41866
rect 33540 41294 33570 41866
rect 33390 41280 33570 41294
rect 33630 41866 33780 41880
rect 33630 41294 33660 41866
rect 33630 41280 33780 41294
rect 34740 41310 34770 42480
rect 34620 41280 34770 41310
rect 34830 41280 34920 42480
rect 34980 41310 35010 42480
rect 34980 41280 35130 41310
rect 35820 42466 35970 42480
rect 35940 41294 35970 42466
rect 35820 41280 35970 41294
rect 36030 42210 36240 42480
rect 36030 41340 36074 42210
rect 36196 41340 36240 42210
rect 36030 41280 36240 41340
rect 36300 41280 36390 42480
rect 36450 42466 36750 42480
rect 36450 41294 36540 42466
rect 36660 41294 36750 42466
rect 36450 41280 36750 41294
rect 36810 41280 36900 42480
rect 36960 42210 37170 42480
rect 36960 41340 37004 42210
rect 37126 41340 37170 42210
rect 36960 41280 37170 41340
rect 37230 42466 37380 42480
rect 37230 41294 37260 42466
rect 38070 42466 38220 42480
rect 37230 41280 37380 41294
rect 37830 41866 37980 41880
rect 37950 41294 37980 41866
rect 37830 41280 37980 41294
rect 38040 41294 38070 41880
rect 38190 41294 38220 42466
rect 38040 41280 38220 41294
rect 38280 41280 38370 42480
rect 38430 42466 38580 42480
rect 38430 41294 38460 42466
rect 38430 41280 38580 41294
rect 39420 42466 39570 42480
rect 39540 41294 39570 42466
rect 39420 41280 39570 41294
rect 39630 42210 39840 42480
rect 39630 41340 39674 42210
rect 39796 41340 39840 42210
rect 39630 41280 39840 41340
rect 39900 41280 39990 42480
rect 40050 42466 40350 42480
rect 40050 41294 40140 42466
rect 40260 41294 40350 42466
rect 40050 41280 40350 41294
rect 40410 41280 40500 42480
rect 40560 42210 40770 42480
rect 40560 41340 40604 42210
rect 40726 41340 40770 42210
rect 40560 41280 40770 41340
rect 40830 42466 40980 42480
rect 40830 41294 40860 42466
rect 43020 42466 43170 42480
rect 40830 41280 40980 41294
rect 41940 41310 41970 41880
rect 41820 41280 41970 41310
rect 42030 41310 42060 41880
rect 42030 41280 42180 41310
rect 43140 41294 43170 42466
rect 43020 41280 43170 41294
rect 43230 41280 43320 42480
rect 43380 42466 43530 42480
rect 43380 41294 43410 42466
rect 44220 42466 44370 42480
rect 43530 41294 43560 41880
rect 43380 41280 43560 41294
rect 43620 41866 43770 41880
rect 43620 41294 43650 41866
rect 43620 41280 43770 41294
rect 44340 41294 44370 42466
rect 44220 41280 44370 41294
rect 44430 41280 44520 42480
rect 44580 42466 44730 42480
rect 44580 41294 44610 42466
rect 45660 42466 45810 42480
rect 44730 41294 44760 41880
rect 44580 41280 44760 41294
rect 44820 41866 44970 41880
rect 44820 41294 44850 41866
rect 44820 41280 44970 41294
rect 45300 41310 45330 41880
rect 45180 41280 45330 41310
rect 45390 41310 45420 41880
rect 45390 41280 45540 41310
rect 45780 41294 45810 42466
rect 45660 41280 45810 41294
rect 45870 42210 46080 42480
rect 45870 41340 45914 42210
rect 46036 41340 46080 42210
rect 45870 41280 46080 41340
rect 46140 41280 46230 42480
rect 46290 42466 46590 42480
rect 46290 41294 46380 42466
rect 46500 41294 46590 42466
rect 46290 41280 46590 41294
rect 46650 41280 46740 42480
rect 46800 42210 47010 42480
rect 46800 41340 46844 42210
rect 46966 41340 47010 42210
rect 46800 41280 47010 41340
rect 47070 42466 47220 42480
rect 47070 41294 47100 42466
rect 47070 41280 47220 41294
rect 47340 42466 47490 42480
rect 47460 41294 47490 42466
rect 47340 41280 47490 41294
rect 47550 42210 47760 42480
rect 47550 41340 47594 42210
rect 47716 41340 47760 42210
rect 47550 41280 47760 41340
rect 47820 41280 47910 42480
rect 47970 42466 48270 42480
rect 47970 41294 48060 42466
rect 48180 41294 48270 42466
rect 47970 41280 48270 41294
rect 48330 41280 48420 42480
rect 48480 42210 48690 42480
rect 48480 41340 48524 42210
rect 48646 41340 48690 42210
rect 48480 41280 48690 41340
rect 48750 42466 48900 42480
rect 48750 41294 48780 42466
rect 48750 41280 48900 41294
rect 5820 40876 5970 40920
rect 5940 39854 5970 40876
rect 5820 39720 5970 39854
rect 6030 39900 6060 40920
rect 6180 39900 6210 40920
rect 6030 39720 6210 39900
rect 6270 40906 6450 40920
rect 6270 39734 6300 40906
rect 6420 39734 6450 40906
rect 6270 39720 6450 39734
rect 6510 40906 6660 40920
rect 6510 39734 6540 40906
rect 8220 40906 8370 40920
rect 8340 40334 8370 40906
rect 8220 40320 8370 40334
rect 8430 40906 8610 40920
rect 8430 40334 8460 40906
rect 8580 40334 8610 40906
rect 8430 40320 8610 40334
rect 8670 40906 8820 40920
rect 8670 40334 8700 40906
rect 8670 40320 8820 40334
rect 9660 40906 9810 40920
rect 9780 40334 9810 40906
rect 9660 40320 9810 40334
rect 9870 40906 10050 40920
rect 9870 40334 9900 40906
rect 10020 40334 10050 40906
rect 9870 40320 10050 40334
rect 10110 40906 10260 40920
rect 10110 40334 10140 40906
rect 10110 40320 10260 40334
rect 10620 40906 10770 40920
rect 6510 39720 6660 39734
rect 10740 39734 10770 40906
rect 10620 39720 10770 39734
rect 10830 40906 11010 40920
rect 10830 39734 10860 40906
rect 10980 39734 11010 40906
rect 10830 39720 11010 39734
rect 11070 39900 11100 40920
rect 11220 39900 11250 40920
rect 11070 39720 11250 39900
rect 11310 40876 11460 40920
rect 11310 39854 11340 40876
rect 11310 39720 11460 39854
rect 11580 40906 11730 40920
rect 11700 39734 11730 40906
rect 11580 39720 11730 39734
rect 11790 40860 12000 40920
rect 11790 39990 11834 40860
rect 11956 39990 12000 40860
rect 11790 39720 12000 39990
rect 12060 39720 12150 40920
rect 12210 40906 12510 40920
rect 12210 39734 12300 40906
rect 12420 39734 12510 40906
rect 12210 39720 12510 39734
rect 12570 39720 12660 40920
rect 12720 40860 12930 40920
rect 12720 39990 12764 40860
rect 12886 39990 12930 40860
rect 12720 39720 12930 39990
rect 12990 40906 13140 40920
rect 12990 39734 13020 40906
rect 13500 40906 13650 40920
rect 13620 40334 13650 40906
rect 13500 40320 13650 40334
rect 13710 40906 13890 40920
rect 13710 40334 13740 40906
rect 13860 40334 13890 40906
rect 13710 40320 13890 40334
rect 13950 40906 14100 40920
rect 13950 40334 13980 40906
rect 13950 40320 14100 40334
rect 14460 40906 14610 40920
rect 14580 40334 14610 40906
rect 14460 40320 14610 40334
rect 14670 40906 14850 40920
rect 14670 40334 14700 40906
rect 14820 40334 14850 40906
rect 14670 40320 14850 40334
rect 14910 40906 15090 40920
rect 14910 40334 14940 40906
rect 15060 40334 15090 40906
rect 14910 40320 15090 40334
rect 15150 40906 15300 40920
rect 15150 40334 15180 40906
rect 15150 40320 15300 40334
rect 15660 40890 15810 40920
rect 15780 40320 15810 40890
rect 15870 40890 16020 40920
rect 15870 40320 15900 40890
rect 16380 40906 16530 40920
rect 12990 39720 13140 39734
rect 16500 39734 16530 40906
rect 16380 39720 16530 39734
rect 16590 39720 16680 40920
rect 16740 40906 16920 40920
rect 16740 39734 16770 40906
rect 16890 40320 16920 40906
rect 16980 40906 17130 40920
rect 16980 40334 17010 40906
rect 16980 40320 17130 40334
rect 17670 40906 17820 40920
rect 17790 40334 17820 40906
rect 17670 40320 17820 40334
rect 17880 40906 18060 40920
rect 17880 40320 17910 40906
rect 16740 39720 16890 39734
rect 18030 39734 18060 40906
rect 17910 39720 18060 39734
rect 18120 39720 18210 40920
rect 18270 40906 18420 40920
rect 18270 39734 18300 40906
rect 18540 40890 18690 40920
rect 18660 40320 18690 40890
rect 18750 40890 18900 40920
rect 18750 40320 18780 40890
rect 19260 40906 19410 40920
rect 18270 39720 18420 39734
rect 19380 39734 19410 40906
rect 19260 39720 19410 39734
rect 19470 39720 19560 40920
rect 19620 40906 19800 40920
rect 19620 39734 19650 40906
rect 19770 40320 19800 40906
rect 19860 40906 20010 40920
rect 19860 40334 19890 40906
rect 19860 40320 20010 40334
rect 20940 40906 21090 40920
rect 21060 40334 21090 40906
rect 20940 40320 21090 40334
rect 21150 40906 21330 40920
rect 21150 40334 21180 40906
rect 21300 40334 21330 40906
rect 21150 40320 21330 40334
rect 21390 40906 21540 40920
rect 21390 40334 21420 40906
rect 21390 40320 21540 40334
rect 21900 40906 22050 40920
rect 19620 39720 19770 39734
rect 22020 39734 22050 40906
rect 21900 39720 22050 39734
rect 22110 40860 22320 40920
rect 22110 39990 22154 40860
rect 22276 39990 22320 40860
rect 22110 39720 22320 39990
rect 22380 39720 22470 40920
rect 22530 40906 22830 40920
rect 22530 39734 22620 40906
rect 22740 39734 22830 40906
rect 22530 39720 22830 39734
rect 22890 39720 22980 40920
rect 23040 40860 23250 40920
rect 23040 39990 23084 40860
rect 23206 39990 23250 40860
rect 23040 39720 23250 39990
rect 23310 40906 23460 40920
rect 23310 39734 23340 40906
rect 23310 39720 23460 39734
rect 23820 40890 23970 40920
rect 23940 39720 23970 40890
rect 24030 39720 24120 40920
rect 24180 40890 24330 40920
rect 24180 39720 24210 40890
rect 24780 40906 24930 40920
rect 24900 39734 24930 40906
rect 24780 39720 24930 39734
rect 24990 39720 25080 40920
rect 25140 40906 25320 40920
rect 25140 39734 25170 40906
rect 25290 40320 25320 40906
rect 25380 40906 25530 40920
rect 25380 40334 25410 40906
rect 25380 40320 25530 40334
rect 26220 40876 26370 40920
rect 25140 39720 25290 39734
rect 26340 39854 26370 40876
rect 26220 39720 26370 39854
rect 26430 39900 26460 40920
rect 26580 39900 26610 40920
rect 26430 39720 26610 39900
rect 26670 40906 26850 40920
rect 26670 39734 26700 40906
rect 26820 39734 26850 40906
rect 26670 39720 26850 39734
rect 26910 40740 27090 40920
rect 26910 39720 26940 40740
rect 27060 39720 27090 40740
rect 27150 40906 27300 40920
rect 27150 39734 27180 40906
rect 27900 40890 28050 40920
rect 28020 40320 28050 40890
rect 28110 40890 28260 40920
rect 28110 40320 28140 40890
rect 30540 40906 30690 40920
rect 30660 40334 30690 40906
rect 30540 40320 30690 40334
rect 30750 40906 30930 40920
rect 30750 40334 30780 40906
rect 30900 40334 30930 40906
rect 30750 40320 30930 40334
rect 30990 40906 31140 40920
rect 30990 40334 31020 40906
rect 30990 40320 31140 40334
rect 31980 40906 32130 40920
rect 32100 40334 32130 40906
rect 31980 40320 32130 40334
rect 32190 40906 32370 40920
rect 32190 40334 32220 40906
rect 32340 40334 32370 40906
rect 32190 40320 32370 40334
rect 32430 40906 32580 40920
rect 32430 40334 32460 40906
rect 32430 40320 32580 40334
rect 33420 40906 33570 40920
rect 27150 39720 27300 39734
rect 33540 39734 33570 40906
rect 33420 39720 33570 39734
rect 33630 40860 33840 40920
rect 33630 39990 33674 40860
rect 33796 39990 33840 40860
rect 33630 39720 33840 39990
rect 33900 39720 33990 40920
rect 34050 40906 34350 40920
rect 34050 39734 34140 40906
rect 34260 39734 34350 40906
rect 34050 39720 34350 39734
rect 34410 39720 34500 40920
rect 34560 40860 34770 40920
rect 34560 39990 34604 40860
rect 34726 39990 34770 40860
rect 34560 39720 34770 39990
rect 34830 40906 34980 40920
rect 34830 39734 34860 40906
rect 34830 39720 34980 39734
rect 36060 40906 36210 40920
rect 36180 39734 36210 40906
rect 36060 39720 36210 39734
rect 36270 39720 36360 40920
rect 36420 40906 36600 40920
rect 36420 39734 36450 40906
rect 36570 40320 36600 40906
rect 36660 40906 36810 40920
rect 36660 40334 36690 40906
rect 36660 40320 36810 40334
rect 37740 40906 37890 40920
rect 37860 40334 37890 40906
rect 37740 40320 37890 40334
rect 37950 40906 38130 40920
rect 37950 40334 37980 40906
rect 38100 40334 38130 40906
rect 37950 40320 38130 40334
rect 38190 40906 38340 40920
rect 38190 40334 38220 40906
rect 38190 40320 38340 40334
rect 38940 40906 39090 40920
rect 36420 39720 36570 39734
rect 39060 39734 39090 40906
rect 38940 39720 39090 39734
rect 39150 39720 39240 40920
rect 39300 40906 39480 40920
rect 39300 39734 39330 40906
rect 39450 40320 39480 40906
rect 39540 40906 39690 40920
rect 39540 40334 39570 40906
rect 39540 40320 39690 40334
rect 40380 40906 40530 40920
rect 40500 40334 40530 40906
rect 40380 40320 40530 40334
rect 40590 40906 40770 40920
rect 40590 40334 40620 40906
rect 40740 40334 40770 40906
rect 40590 40320 40770 40334
rect 40830 40906 40980 40920
rect 40830 40334 40860 40906
rect 40830 40320 40980 40334
rect 41820 40890 41970 40920
rect 41940 40320 41970 40890
rect 42030 40890 42180 40920
rect 42030 40320 42060 40890
rect 43020 40906 43170 40920
rect 39300 39720 39450 39734
rect 43140 39734 43170 40906
rect 43020 39720 43170 39734
rect 43230 39720 43320 40920
rect 43380 40906 43560 40920
rect 43380 39734 43410 40906
rect 43530 40320 43560 40906
rect 43620 40906 43770 40920
rect 43620 40334 43650 40906
rect 43620 40320 43770 40334
rect 44700 40890 44850 40920
rect 44820 40320 44850 40890
rect 44910 40890 45060 40920
rect 44910 40320 44940 40890
rect 45990 40906 46140 40920
rect 46110 40334 46140 40906
rect 45990 40320 46140 40334
rect 46200 40906 46380 40920
rect 46200 40320 46230 40906
rect 43380 39720 43530 39734
rect 46350 39734 46380 40906
rect 46230 39720 46380 39734
rect 46440 39720 46530 40920
rect 46590 40906 46740 40920
rect 46590 39734 46620 40906
rect 46590 39720 46740 39734
rect 47580 40906 47730 40920
rect 47700 39734 47730 40906
rect 47580 39720 47730 39734
rect 47790 39720 47880 40920
rect 47940 40906 48120 40920
rect 47940 39734 47970 40906
rect 48090 40320 48120 40906
rect 48180 40906 48330 40920
rect 48180 40334 48210 40906
rect 48180 40320 48330 40334
rect 49260 40906 49410 40920
rect 49380 40334 49410 40906
rect 49260 40320 49410 40334
rect 49470 40906 49650 40920
rect 49470 40334 49500 40906
rect 49620 40334 49650 40906
rect 49470 40320 49650 40334
rect 49710 40906 49860 40920
rect 49710 40334 49740 40906
rect 49710 40320 49860 40334
rect 47940 39720 48090 39734
rect 8550 36466 8700 36480
rect 5580 35866 5730 35880
rect 5700 35294 5730 35866
rect 5580 35280 5730 35294
rect 5790 35866 5970 35880
rect 5790 35294 5820 35866
rect 5940 35294 5970 35866
rect 5790 35280 5970 35294
rect 6030 35866 6180 35880
rect 6030 35294 6060 35866
rect 6030 35280 6180 35294
rect 7140 35310 7170 35880
rect 7020 35280 7170 35310
rect 7230 35310 7260 35880
rect 7230 35280 7380 35310
rect 8310 35866 8460 35880
rect 8430 35294 8460 35866
rect 8310 35280 8460 35294
rect 8520 35294 8550 35880
rect 8670 35294 8700 36466
rect 8520 35280 8700 35294
rect 8760 35280 8850 36480
rect 8910 36466 9060 36480
rect 8910 35294 8940 36466
rect 12390 36466 12540 36480
rect 8910 35280 9060 35294
rect 10860 35866 11010 35880
rect 10980 35294 11010 35866
rect 10860 35280 11010 35294
rect 11070 35866 11250 35880
rect 11070 35294 11100 35866
rect 11220 35294 11250 35866
rect 11070 35280 11250 35294
rect 11310 35866 11460 35880
rect 11310 35294 11340 35866
rect 11310 35280 11460 35294
rect 12150 35866 12300 35880
rect 12270 35294 12300 35866
rect 12150 35280 12300 35294
rect 12360 35294 12390 35880
rect 12510 35294 12540 36466
rect 12360 35280 12540 35294
rect 12600 35280 12690 36480
rect 12750 36466 12900 36480
rect 12750 35294 12780 36466
rect 15270 36466 15420 36480
rect 12750 35280 12900 35294
rect 15030 35866 15180 35880
rect 15150 35294 15180 35866
rect 15030 35280 15180 35294
rect 15240 35294 15270 35880
rect 15390 35294 15420 36466
rect 15240 35280 15420 35294
rect 15480 35280 15570 36480
rect 15630 36466 15780 36480
rect 15630 35294 15660 36466
rect 26460 36466 26610 36480
rect 15630 35280 15780 35294
rect 16620 35866 16770 35880
rect 16740 35294 16770 35866
rect 16620 35280 16770 35294
rect 16830 35866 17010 35880
rect 16830 35294 16860 35866
rect 16980 35294 17010 35866
rect 16830 35280 17010 35294
rect 17070 35866 17250 35880
rect 17070 35294 17100 35866
rect 17220 35294 17250 35866
rect 17070 35280 17250 35294
rect 17310 35866 17460 35880
rect 17310 35294 17340 35866
rect 17310 35280 17460 35294
rect 18060 35866 18210 35880
rect 18180 35294 18210 35866
rect 18060 35280 18210 35294
rect 18270 35866 18450 35880
rect 18270 35294 18300 35866
rect 18420 35294 18450 35866
rect 18270 35280 18450 35294
rect 18510 35866 18660 35880
rect 18510 35294 18540 35866
rect 18510 35280 18660 35294
rect 19500 35866 19650 35880
rect 19620 35294 19650 35866
rect 19500 35280 19650 35294
rect 19710 35866 19890 35880
rect 19710 35294 19740 35866
rect 19860 35294 19890 35866
rect 19710 35280 19890 35294
rect 19950 35866 20100 35880
rect 19950 35294 19980 35866
rect 19950 35280 20100 35294
rect 20940 35866 21090 35880
rect 21060 35294 21090 35866
rect 20940 35280 21090 35294
rect 21150 35866 21330 35880
rect 21150 35294 21180 35866
rect 21300 35294 21330 35866
rect 21150 35280 21330 35294
rect 21390 35866 21540 35880
rect 21390 35294 21420 35866
rect 21390 35280 21540 35294
rect 22380 35866 22530 35880
rect 22500 35294 22530 35866
rect 22380 35280 22530 35294
rect 22590 35866 22770 35880
rect 22590 35294 22620 35866
rect 22740 35294 22770 35866
rect 22590 35280 22770 35294
rect 22830 35866 22980 35880
rect 22830 35294 22860 35866
rect 22830 35280 22980 35294
rect 23940 35310 23970 35880
rect 23820 35280 23970 35310
rect 24030 35310 24060 35880
rect 24030 35280 24180 35310
rect 25020 35866 25170 35880
rect 25140 35294 25170 35866
rect 25020 35280 25170 35294
rect 25230 35866 25410 35880
rect 25230 35294 25260 35866
rect 25380 35294 25410 35866
rect 25230 35280 25410 35294
rect 25470 35866 25620 35880
rect 25470 35294 25500 35866
rect 25470 35280 25620 35294
rect 26580 35294 26610 36466
rect 26460 35280 26610 35294
rect 26670 35280 26760 36480
rect 26820 36466 26970 36480
rect 26820 35294 26850 36466
rect 30060 36466 30210 36480
rect 26970 35294 27000 35880
rect 26820 35280 27000 35294
rect 27060 35866 27210 35880
rect 27060 35294 27090 35866
rect 27060 35280 27210 35294
rect 27900 35866 28050 35880
rect 28020 35294 28050 35866
rect 27900 35280 28050 35294
rect 28110 35866 28290 35880
rect 28110 35294 28140 35866
rect 28260 35294 28290 35866
rect 28110 35280 28290 35294
rect 28350 35866 28500 35880
rect 28350 35294 28380 35866
rect 28350 35280 28500 35294
rect 29100 35866 29250 35880
rect 29220 35294 29250 35866
rect 29100 35280 29250 35294
rect 29310 35866 29490 35880
rect 29310 35294 29340 35866
rect 29460 35294 29490 35866
rect 29310 35280 29490 35294
rect 29550 35866 29700 35880
rect 29550 35294 29580 35866
rect 29550 35280 29700 35294
rect 30180 35294 30210 36466
rect 30060 35280 30210 35294
rect 30270 35280 30360 36480
rect 30420 36466 30570 36480
rect 30420 35294 30450 36466
rect 32310 36466 32460 36480
rect 30570 35294 30600 35880
rect 30420 35280 30600 35294
rect 30660 35866 30810 35880
rect 30660 35294 30690 35866
rect 30660 35280 30810 35294
rect 31380 35310 31410 35880
rect 31260 35280 31410 35310
rect 31470 35310 31500 35880
rect 31470 35280 31620 35310
rect 32070 35866 32220 35880
rect 32190 35294 32220 35866
rect 32070 35280 32220 35294
rect 32280 35294 32310 35880
rect 32430 35294 32460 36466
rect 32280 35280 32460 35294
rect 32520 35280 32610 36480
rect 32670 36466 32820 36480
rect 32670 35294 32700 36466
rect 35580 36466 35730 36480
rect 32670 35280 32820 35294
rect 33180 35866 33330 35880
rect 33300 35294 33330 35866
rect 33180 35280 33330 35294
rect 33390 35866 33570 35880
rect 33390 35294 33420 35866
rect 33540 35294 33570 35866
rect 33390 35280 33570 35294
rect 33630 35866 33780 35880
rect 33630 35294 33660 35866
rect 33630 35280 33780 35294
rect 34620 35866 34770 35880
rect 34740 35294 34770 35866
rect 34620 35280 34770 35294
rect 34830 35866 35010 35880
rect 34830 35294 34860 35866
rect 34980 35294 35010 35866
rect 34830 35280 35010 35294
rect 35070 35866 35220 35880
rect 35070 35294 35100 35866
rect 35070 35280 35220 35294
rect 35700 35294 35730 36466
rect 35580 35280 35730 35294
rect 35790 36210 36000 36480
rect 35790 35340 35834 36210
rect 35956 35340 36000 36210
rect 35790 35280 36000 35340
rect 36060 35280 36150 36480
rect 36210 36466 36510 36480
rect 36210 35294 36300 36466
rect 36420 35294 36510 36466
rect 36210 35280 36510 35294
rect 36570 35280 36660 36480
rect 36720 36210 36930 36480
rect 36720 35340 36764 36210
rect 36886 35340 36930 36210
rect 36720 35280 36930 35340
rect 36990 36466 37140 36480
rect 36990 35294 37020 36466
rect 39900 36466 40050 36480
rect 36990 35280 37140 35294
rect 39060 35310 39090 35880
rect 38940 35280 39090 35310
rect 39150 35310 39180 35880
rect 39150 35280 39300 35310
rect 40020 35294 40050 36466
rect 39900 35280 40050 35294
rect 40110 35460 40140 36480
rect 40260 35460 40290 36480
rect 40110 35280 40290 35460
rect 40350 36466 40530 36480
rect 40350 35294 40380 36466
rect 40500 35294 40530 36466
rect 40350 35280 40530 35294
rect 40590 36300 40770 36480
rect 40590 35280 40620 36300
rect 40740 35280 40770 36300
rect 40830 36346 40980 36480
rect 40830 35324 40860 36346
rect 42630 36466 42780 36480
rect 40830 35280 40980 35324
rect 41700 35310 41730 35880
rect 41580 35280 41730 35310
rect 41790 35310 41820 35880
rect 41790 35280 41940 35310
rect 42390 35866 42540 35880
rect 42510 35294 42540 35866
rect 42390 35280 42540 35294
rect 42600 35294 42630 35880
rect 42750 35294 42780 36466
rect 42600 35280 42780 35294
rect 42840 35280 42930 36480
rect 42990 36466 43140 36480
rect 42990 35294 43020 36466
rect 44460 36466 44610 36480
rect 42990 35280 43140 35294
rect 43620 35310 43650 35880
rect 43500 35280 43650 35310
rect 43710 35310 43740 35880
rect 43710 35280 43860 35310
rect 44580 35294 44610 36466
rect 44460 35280 44610 35294
rect 44670 35280 44760 36480
rect 44820 36466 44970 36480
rect 44820 35294 44850 36466
rect 47580 36466 47730 36480
rect 44970 35294 45000 35880
rect 44820 35280 45000 35294
rect 45060 35866 45210 35880
rect 45060 35294 45090 35866
rect 45060 35280 45210 35294
rect 46140 35866 46290 35880
rect 46260 35294 46290 35866
rect 46140 35280 46290 35294
rect 46350 35866 46530 35880
rect 46350 35294 46380 35866
rect 46500 35294 46530 35866
rect 46350 35280 46530 35294
rect 46590 35866 46740 35880
rect 46590 35294 46620 35866
rect 46590 35280 46740 35294
rect 47700 35294 47730 36466
rect 47580 35280 47730 35294
rect 47790 35280 47880 36480
rect 47940 36466 48090 36480
rect 47940 35294 47970 36466
rect 48090 35294 48120 35880
rect 47940 35280 48120 35294
rect 48180 35866 48330 35880
rect 48180 35294 48210 35866
rect 48180 35280 48330 35294
rect 49260 35866 49410 35880
rect 49380 35294 49410 35866
rect 49260 35280 49410 35294
rect 49470 35866 49650 35880
rect 49470 35294 49500 35866
rect 49620 35294 49650 35866
rect 49470 35280 49650 35294
rect 49710 35866 49860 35880
rect 49710 35294 49740 35866
rect 49710 35280 49860 35294
rect 6630 34906 6780 34920
rect 6750 34334 6780 34906
rect 6630 34320 6780 34334
rect 6840 34906 7020 34920
rect 6840 34320 6870 34906
rect 6990 33734 7020 34906
rect 6870 33720 7020 33734
rect 7080 33720 7170 34920
rect 7230 34906 7380 34920
rect 7230 33734 7260 34906
rect 7830 34906 7980 34920
rect 7950 34334 7980 34906
rect 7830 34320 7980 34334
rect 8040 34906 8220 34920
rect 8040 34320 8070 34906
rect 7230 33720 7380 33734
rect 8190 33734 8220 34906
rect 8070 33720 8220 33734
rect 8280 33720 8370 34920
rect 8430 34906 8580 34920
rect 8430 33734 8460 34906
rect 8430 33720 8580 33734
rect 8940 34906 9090 34920
rect 9060 33734 9090 34906
rect 8940 33720 9090 33734
rect 9150 34860 9360 34920
rect 9150 33990 9194 34860
rect 9316 33990 9360 34860
rect 9150 33720 9360 33990
rect 9420 33720 9510 34920
rect 9570 34906 9870 34920
rect 9570 33734 9660 34906
rect 9780 33734 9870 34906
rect 9570 33720 9870 33734
rect 9930 33720 10020 34920
rect 10080 34860 10290 34920
rect 10080 33990 10124 34860
rect 10246 33990 10290 34860
rect 10080 33720 10290 33990
rect 10350 34906 10500 34920
rect 10350 33734 10380 34906
rect 10350 33720 10500 33734
rect 11100 34906 11250 34920
rect 11220 33734 11250 34906
rect 11100 33720 11250 33734
rect 11310 34860 11520 34920
rect 11310 33990 11354 34860
rect 11476 33990 11520 34860
rect 11310 33720 11520 33990
rect 11580 33720 11670 34920
rect 11730 34906 12030 34920
rect 11730 33734 11820 34906
rect 11940 33734 12030 34906
rect 11730 33720 12030 33734
rect 12090 33720 12180 34920
rect 12240 34860 12450 34920
rect 12240 33990 12284 34860
rect 12406 33990 12450 34860
rect 12240 33720 12450 33990
rect 12510 34906 12660 34920
rect 12510 33734 12540 34906
rect 13740 34890 13890 34920
rect 13860 34320 13890 34890
rect 13950 34890 14100 34920
rect 13950 34320 13980 34890
rect 15180 34906 15330 34920
rect 15300 34334 15330 34906
rect 15180 34320 15330 34334
rect 15390 34906 15570 34920
rect 15390 34334 15420 34906
rect 15540 34334 15570 34906
rect 15390 34320 15570 34334
rect 15630 34906 15780 34920
rect 15630 34334 15660 34906
rect 15630 34320 15780 34334
rect 16620 34906 16770 34920
rect 12510 33720 12660 33734
rect 16740 33734 16770 34906
rect 16620 33720 16770 33734
rect 16830 33720 16920 34920
rect 16980 34906 17160 34920
rect 16980 33734 17010 34906
rect 17130 34320 17160 34906
rect 17220 34906 17370 34920
rect 17220 34334 17250 34906
rect 17220 34320 17370 34334
rect 19260 34906 19410 34920
rect 19380 34334 19410 34906
rect 19260 34320 19410 34334
rect 19470 34906 19650 34920
rect 19470 34334 19500 34906
rect 19620 34334 19650 34906
rect 19470 34320 19650 34334
rect 19710 34906 19860 34920
rect 19710 34334 19740 34906
rect 19710 34320 19860 34334
rect 20700 34906 20850 34920
rect 20820 34334 20850 34906
rect 20700 34320 20850 34334
rect 20910 34906 21090 34920
rect 20910 34334 20940 34906
rect 21060 34334 21090 34906
rect 20910 34320 21090 34334
rect 21150 34906 21330 34920
rect 21150 34334 21180 34906
rect 21300 34334 21330 34906
rect 21150 34320 21330 34334
rect 21390 34906 21540 34920
rect 21390 34334 21420 34906
rect 21390 34320 21540 34334
rect 23340 34906 23490 34920
rect 16980 33720 17130 33734
rect 23460 33734 23490 34906
rect 23340 33720 23490 33734
rect 23550 33720 23640 34920
rect 23700 34906 23880 34920
rect 23700 33734 23730 34906
rect 23850 34320 23880 34906
rect 23940 34906 24090 34920
rect 23940 34334 23970 34906
rect 23940 34320 24090 34334
rect 24780 34906 24930 34920
rect 23700 33720 23850 33734
rect 24900 33734 24930 34906
rect 24780 33720 24930 33734
rect 24990 33720 25080 34920
rect 25140 34906 25320 34920
rect 25140 33734 25170 34906
rect 25290 34320 25320 34906
rect 25380 34906 25530 34920
rect 25380 34334 25410 34906
rect 25380 34320 25530 34334
rect 25980 34906 26130 34920
rect 25140 33720 25290 33734
rect 26100 33734 26130 34906
rect 25980 33720 26130 33734
rect 26190 34860 26400 34920
rect 26190 33990 26234 34860
rect 26356 33990 26400 34860
rect 26190 33720 26400 33990
rect 26460 33720 26550 34920
rect 26610 34906 26910 34920
rect 26610 33734 26700 34906
rect 26820 33734 26910 34906
rect 26610 33720 26910 33734
rect 26970 33720 27060 34920
rect 27120 34860 27330 34920
rect 27120 33990 27164 34860
rect 27286 33990 27330 34860
rect 27120 33720 27330 33990
rect 27390 34906 27540 34920
rect 27390 33734 27420 34906
rect 30300 34890 30450 34920
rect 30420 34320 30450 34890
rect 30510 34890 30660 34920
rect 30510 34320 30540 34890
rect 31020 34906 31170 34920
rect 31140 34334 31170 34906
rect 31020 34320 31170 34334
rect 31230 34906 31410 34920
rect 31230 34334 31260 34906
rect 31380 34334 31410 34906
rect 31230 34320 31410 34334
rect 31470 34906 31620 34920
rect 31470 34334 31500 34906
rect 31470 34320 31620 34334
rect 31980 34906 32130 34920
rect 27390 33720 27540 33734
rect 32100 33734 32130 34906
rect 31980 33720 32130 33734
rect 32190 33720 32280 34920
rect 32340 34906 32520 34920
rect 32340 33734 32370 34906
rect 32490 34320 32520 34906
rect 32580 34906 32730 34920
rect 32580 34334 32610 34906
rect 32580 34320 32730 34334
rect 33180 34906 33330 34920
rect 33300 34334 33330 34906
rect 33180 34320 33330 34334
rect 33390 34906 33570 34920
rect 33390 34334 33420 34906
rect 33540 34334 33570 34906
rect 33390 34320 33570 34334
rect 33630 34906 33780 34920
rect 33630 34334 33660 34906
rect 33630 34320 33780 34334
rect 34620 34906 34770 34920
rect 34740 34334 34770 34906
rect 34620 34320 34770 34334
rect 34830 34906 35010 34920
rect 34830 34334 34860 34906
rect 34980 34334 35010 34906
rect 34830 34320 35010 34334
rect 35070 34906 35220 34920
rect 35070 34334 35100 34906
rect 35070 34320 35220 34334
rect 36060 34906 36210 34920
rect 36180 34334 36210 34906
rect 36060 34320 36210 34334
rect 36270 34906 36450 34920
rect 36270 34334 36300 34906
rect 36420 34334 36450 34906
rect 36270 34320 36450 34334
rect 36510 34906 36660 34920
rect 36510 34334 36540 34906
rect 36510 34320 36660 34334
rect 37500 34906 37650 34920
rect 37620 34334 37650 34906
rect 37500 34320 37650 34334
rect 37710 34906 37890 34920
rect 37710 34334 37740 34906
rect 37860 34334 37890 34906
rect 37710 34320 37890 34334
rect 37950 34906 38100 34920
rect 37950 34334 37980 34906
rect 37950 34320 38100 34334
rect 38940 34906 39090 34920
rect 39060 34334 39090 34906
rect 38940 34320 39090 34334
rect 39150 34906 39330 34920
rect 39150 34334 39180 34906
rect 39300 34334 39330 34906
rect 39150 34320 39330 34334
rect 39390 34906 39540 34920
rect 39390 34334 39420 34906
rect 39390 34320 39540 34334
rect 40140 34906 40290 34920
rect 32340 33720 32490 33734
rect 40260 33734 40290 34906
rect 40140 33720 40290 33734
rect 40350 33720 40440 34920
rect 40500 34906 40680 34920
rect 40500 33734 40530 34906
rect 40650 34320 40680 34906
rect 40740 34906 40890 34920
rect 40740 34334 40770 34906
rect 40740 34320 40890 34334
rect 41580 34906 41730 34920
rect 41700 34334 41730 34906
rect 41580 34320 41730 34334
rect 41790 34906 41970 34920
rect 41790 34334 41820 34906
rect 41940 34334 41970 34906
rect 41790 34320 41970 34334
rect 42030 34906 42180 34920
rect 42030 34334 42060 34906
rect 42030 34320 42180 34334
rect 43020 34906 43170 34920
rect 40500 33720 40650 33734
rect 43140 33734 43170 34906
rect 43020 33720 43170 33734
rect 43230 33720 43320 34920
rect 43380 34906 43560 34920
rect 43380 33734 43410 34906
rect 43530 34320 43560 34906
rect 43620 34906 43770 34920
rect 43620 34334 43650 34906
rect 43620 34320 43770 34334
rect 44220 34906 44370 34920
rect 43380 33720 43530 33734
rect 44340 33734 44370 34906
rect 44220 33720 44370 33734
rect 44430 34860 44640 34920
rect 44430 33990 44474 34860
rect 44596 33990 44640 34860
rect 44430 33720 44640 33990
rect 44700 33720 44790 34920
rect 44850 34906 45150 34920
rect 44850 33734 44940 34906
rect 45060 33734 45150 34906
rect 44850 33720 45150 33734
rect 45210 33720 45300 34920
rect 45360 34860 45570 34920
rect 45360 33990 45404 34860
rect 45526 33990 45570 34860
rect 45360 33720 45570 33990
rect 45630 34906 45780 34920
rect 45630 33734 45660 34906
rect 45630 33720 45780 33734
rect 46140 34906 46290 34920
rect 46260 33734 46290 34906
rect 46140 33720 46290 33734
rect 46350 33720 46440 34920
rect 46500 34906 46680 34920
rect 46500 33734 46530 34906
rect 46650 34320 46680 34906
rect 46740 34906 46890 34920
rect 46740 34334 46770 34906
rect 46740 34320 46890 34334
rect 47580 34906 47730 34920
rect 47700 34334 47730 34906
rect 47580 34320 47730 34334
rect 47790 34906 47970 34920
rect 47790 34334 47820 34906
rect 47940 34334 47970 34906
rect 47790 34320 47970 34334
rect 48030 34906 48180 34920
rect 48030 34334 48060 34906
rect 48030 34320 48180 34334
rect 49020 34906 49170 34920
rect 49140 34334 49170 34906
rect 49020 34320 49170 34334
rect 49230 34906 49410 34920
rect 49230 34334 49260 34906
rect 49380 34334 49410 34906
rect 49230 34320 49410 34334
rect 49470 34906 49620 34920
rect 49470 34334 49500 34906
rect 49470 34320 49620 34334
rect 46500 33720 46650 33734
rect 5340 30466 5490 30480
rect 5460 29294 5490 30466
rect 5340 29280 5490 29294
rect 5550 30210 5760 30480
rect 5550 29340 5594 30210
rect 5716 29340 5760 30210
rect 5550 29280 5760 29340
rect 5820 29280 5910 30480
rect 5970 30466 6270 30480
rect 5970 29294 6060 30466
rect 6180 29294 6270 30466
rect 5970 29280 6270 29294
rect 6330 29280 6420 30480
rect 6480 30210 6690 30480
rect 6480 29340 6524 30210
rect 6646 29340 6690 30210
rect 6480 29280 6690 29340
rect 6750 30466 6900 30480
rect 6750 29294 6780 30466
rect 6750 29280 6900 29294
rect 7980 30466 8130 30480
rect 8100 29294 8130 30466
rect 7980 29280 8130 29294
rect 8190 29280 8280 30480
rect 8340 30466 8490 30480
rect 8340 29294 8370 30466
rect 11100 30466 11250 30480
rect 8490 29294 8520 29880
rect 8340 29280 8520 29294
rect 8580 29866 8730 29880
rect 8580 29294 8610 29866
rect 8580 29280 8730 29294
rect 9660 29866 9810 29880
rect 9780 29294 9810 29866
rect 9660 29280 9810 29294
rect 9870 29866 10050 29880
rect 9870 29294 9900 29866
rect 10020 29294 10050 29866
rect 9870 29280 10050 29294
rect 10110 29866 10260 29880
rect 10110 29294 10140 29866
rect 10110 29280 10260 29294
rect 11220 29294 11250 30466
rect 11100 29280 11250 29294
rect 11310 30210 11520 30480
rect 11310 29340 11354 30210
rect 11476 29340 11520 30210
rect 11310 29280 11520 29340
rect 11580 29280 11670 30480
rect 11730 30466 12030 30480
rect 11730 29294 11820 30466
rect 11940 29294 12030 30466
rect 11730 29280 12030 29294
rect 12090 29280 12180 30480
rect 12240 30210 12450 30480
rect 12240 29340 12284 30210
rect 12406 29340 12450 30210
rect 12240 29280 12450 29340
rect 12510 30466 12660 30480
rect 12510 29294 12540 30466
rect 12510 29280 12660 29294
rect 14700 30466 14850 30480
rect 14820 29294 14850 30466
rect 14700 29280 14850 29294
rect 14910 30210 15120 30480
rect 14910 29340 14954 30210
rect 15076 29340 15120 30210
rect 14910 29280 15120 29340
rect 15180 29280 15270 30480
rect 15330 30466 15630 30480
rect 15330 29294 15420 30466
rect 15540 29294 15630 30466
rect 15330 29280 15630 29294
rect 15690 29280 15780 30480
rect 15840 30210 16050 30480
rect 15840 29340 15884 30210
rect 16006 29340 16050 30210
rect 15840 29280 16050 29340
rect 16110 30466 16260 30480
rect 16110 29294 16140 30466
rect 16110 29280 16260 29294
rect 17100 30466 17250 30480
rect 17220 29294 17250 30466
rect 17100 29280 17250 29294
rect 17310 30210 17520 30480
rect 17310 29340 17354 30210
rect 17476 29340 17520 30210
rect 17310 29280 17520 29340
rect 17580 29280 17670 30480
rect 17730 30466 18030 30480
rect 17730 29294 17820 30466
rect 17940 29294 18030 30466
rect 17730 29280 18030 29294
rect 18090 29280 18180 30480
rect 18240 30210 18450 30480
rect 18240 29340 18284 30210
rect 18406 29340 18450 30210
rect 18240 29280 18450 29340
rect 18510 30466 18660 30480
rect 18510 29294 18540 30466
rect 18510 29280 18660 29294
rect 19260 30466 19410 30480
rect 19380 29294 19410 30466
rect 19260 29280 19410 29294
rect 19470 30210 19680 30480
rect 19470 29340 19514 30210
rect 19636 29340 19680 30210
rect 19470 29280 19680 29340
rect 19740 29280 19830 30480
rect 19890 30466 20190 30480
rect 19890 29294 19980 30466
rect 20100 29294 20190 30466
rect 19890 29280 20190 29294
rect 20250 29280 20340 30480
rect 20400 30210 20610 30480
rect 20400 29340 20444 30210
rect 20566 29340 20610 30210
rect 20400 29280 20610 29340
rect 20670 30466 20820 30480
rect 20670 29294 20700 30466
rect 22470 30466 22620 30480
rect 20670 29280 20820 29294
rect 21180 29866 21330 29880
rect 21300 29294 21330 29866
rect 21180 29280 21330 29294
rect 21390 29866 21570 29880
rect 21390 29294 21420 29866
rect 21540 29294 21570 29866
rect 21390 29280 21570 29294
rect 21630 29866 21780 29880
rect 21630 29294 21660 29866
rect 21630 29280 21780 29294
rect 22230 29866 22380 29880
rect 22350 29294 22380 29866
rect 22230 29280 22380 29294
rect 22440 29294 22470 29880
rect 22590 29294 22620 30466
rect 22440 29280 22620 29294
rect 22680 29280 22770 30480
rect 22830 30466 22980 30480
rect 22830 29294 22860 30466
rect 26310 30466 26460 30480
rect 22830 29280 22980 29294
rect 23940 29310 23970 29880
rect 23820 29280 23970 29310
rect 24030 29310 24060 29880
rect 24030 29280 24180 29310
rect 24780 29866 24930 29880
rect 24900 29294 24930 29866
rect 24780 29280 24930 29294
rect 24990 29866 25170 29880
rect 24990 29294 25020 29866
rect 25140 29294 25170 29866
rect 24990 29280 25170 29294
rect 25230 29866 25410 29880
rect 25230 29294 25260 29866
rect 25380 29294 25410 29866
rect 25230 29280 25410 29294
rect 25470 29866 25620 29880
rect 25470 29294 25500 29866
rect 25470 29280 25620 29294
rect 26070 29866 26220 29880
rect 26190 29294 26220 29866
rect 26070 29280 26220 29294
rect 26280 29294 26310 29880
rect 26430 29294 26460 30466
rect 26280 29280 26460 29294
rect 26520 29280 26610 30480
rect 26670 30466 26820 30480
rect 26670 29294 26700 30466
rect 29430 30466 29580 30480
rect 26670 29280 26820 29294
rect 27300 29310 27330 29880
rect 27180 29280 27330 29310
rect 27390 29310 27420 29880
rect 27390 29280 27540 29310
rect 27660 29866 27810 29880
rect 27780 29294 27810 29866
rect 27660 29280 27810 29294
rect 27870 29866 28050 29880
rect 27870 29294 27900 29866
rect 28020 29294 28050 29866
rect 27870 29280 28050 29294
rect 28110 29866 28260 29880
rect 28110 29294 28140 29866
rect 28110 29280 28260 29294
rect 28740 29310 28770 29880
rect 28620 29280 28770 29310
rect 28830 29310 28860 29880
rect 28830 29280 28980 29310
rect 29190 29866 29340 29880
rect 29310 29294 29340 29866
rect 29190 29280 29340 29294
rect 29400 29294 29430 29880
rect 29550 29294 29580 30466
rect 29400 29280 29580 29294
rect 29640 29280 29730 30480
rect 29790 30466 29940 30480
rect 29790 29294 29820 30466
rect 29790 29280 29940 29294
rect 30780 30466 30930 30480
rect 30900 29294 30930 30466
rect 30780 29280 30930 29294
rect 30990 30210 31200 30480
rect 30990 29340 31034 30210
rect 31156 29340 31200 30210
rect 30990 29280 31200 29340
rect 31260 29280 31350 30480
rect 31410 30466 31710 30480
rect 31410 29294 31500 30466
rect 31620 29294 31710 30466
rect 31410 29280 31710 29294
rect 31770 29280 31860 30480
rect 31920 30210 32130 30480
rect 31920 29340 31964 30210
rect 32086 29340 32130 30210
rect 31920 29280 32130 29340
rect 32190 30466 32340 30480
rect 32190 29294 32220 30466
rect 36390 30466 36540 30480
rect 32190 29280 32340 29294
rect 33180 29866 33330 29880
rect 33300 29294 33330 29866
rect 33180 29280 33330 29294
rect 33390 29866 33570 29880
rect 33390 29294 33420 29866
rect 33540 29294 33570 29866
rect 33390 29280 33570 29294
rect 33630 29866 33780 29880
rect 33630 29294 33660 29866
rect 33630 29280 33780 29294
rect 34620 29866 34770 29880
rect 34740 29294 34770 29866
rect 34620 29280 34770 29294
rect 34830 29866 35010 29880
rect 34830 29294 34860 29866
rect 34980 29294 35010 29866
rect 34830 29280 35010 29294
rect 35070 29866 35220 29880
rect 35070 29294 35100 29866
rect 35070 29280 35220 29294
rect 36150 29866 36300 29880
rect 36270 29294 36300 29866
rect 36150 29280 36300 29294
rect 36360 29294 36390 29880
rect 36510 29294 36540 30466
rect 36360 29280 36540 29294
rect 36600 29280 36690 30480
rect 36750 30466 36900 30480
rect 36750 29294 36780 30466
rect 38940 30466 39090 30480
rect 36750 29280 36900 29294
rect 37740 29866 37890 29880
rect 37860 29294 37890 29866
rect 37740 29280 37890 29294
rect 37950 29866 38130 29880
rect 37950 29294 37980 29866
rect 38100 29294 38130 29866
rect 37950 29280 38130 29294
rect 38190 29866 38340 29880
rect 38190 29294 38220 29866
rect 38190 29280 38340 29294
rect 39060 29294 39090 30466
rect 38940 29280 39090 29294
rect 39150 29280 39240 30480
rect 39300 30466 39450 30480
rect 39300 29294 39330 30466
rect 43350 30466 43500 30480
rect 39450 29294 39480 29880
rect 39300 29280 39480 29294
rect 39540 29866 39690 29880
rect 39540 29294 39570 29866
rect 39540 29280 39690 29294
rect 40740 29310 40770 29880
rect 40620 29280 40770 29310
rect 40830 29310 40860 29880
rect 40830 29280 40980 29310
rect 41580 29866 41730 29880
rect 41700 29294 41730 29866
rect 41580 29280 41730 29294
rect 41790 29866 41970 29880
rect 41790 29294 41820 29866
rect 41940 29294 41970 29866
rect 41790 29280 41970 29294
rect 42030 29866 42180 29880
rect 42030 29294 42060 29866
rect 42030 29280 42180 29294
rect 43110 29866 43260 29880
rect 43230 29294 43260 29866
rect 43110 29280 43260 29294
rect 43320 29294 43350 29880
rect 43470 29294 43500 30466
rect 43320 29280 43500 29294
rect 43560 29280 43650 30480
rect 43710 30466 43860 30480
rect 43710 29294 43740 30466
rect 43710 29280 43860 29294
rect 44460 30466 44610 30480
rect 44580 29294 44610 30466
rect 44460 29280 44610 29294
rect 44670 29280 44760 30480
rect 44820 30466 44970 30480
rect 44820 29294 44850 30466
rect 48060 30466 48210 30480
rect 44970 29294 45000 29880
rect 44820 29280 45000 29294
rect 45060 29866 45210 29880
rect 45060 29294 45090 29866
rect 45060 29280 45210 29294
rect 46140 29866 46290 29880
rect 46260 29294 46290 29866
rect 46140 29280 46290 29294
rect 46350 29866 46530 29880
rect 46350 29294 46380 29866
rect 46500 29294 46530 29866
rect 46350 29280 46530 29294
rect 46590 29866 46740 29880
rect 46590 29294 46620 29866
rect 46590 29280 46740 29294
rect 48180 29294 48210 30466
rect 48060 29280 48210 29294
rect 48270 30210 48480 30480
rect 48270 29340 48314 30210
rect 48436 29340 48480 30210
rect 48270 29280 48480 29340
rect 48540 29280 48630 30480
rect 48690 30466 48990 30480
rect 48690 29294 48780 30466
rect 48900 29294 48990 30466
rect 48690 29280 48990 29294
rect 49050 29280 49140 30480
rect 49200 30210 49410 30480
rect 49200 29340 49244 30210
rect 49366 29340 49410 30210
rect 49200 29280 49410 29340
rect 49470 30466 49620 30480
rect 49470 29294 49500 30466
rect 49470 29280 49620 29294
rect 7020 28906 7170 28920
rect 7140 27734 7170 28906
rect 7020 27720 7170 27734
rect 7230 28860 7440 28920
rect 7230 27990 7274 28860
rect 7396 27990 7440 28860
rect 7230 27720 7440 27990
rect 7500 27720 7590 28920
rect 7650 28906 7950 28920
rect 7650 27734 7740 28906
rect 7860 27734 7950 28906
rect 7650 27720 7950 27734
rect 8010 27720 8100 28920
rect 8160 28860 8370 28920
rect 8160 27990 8204 28860
rect 8326 27990 8370 28860
rect 8160 27720 8370 27990
rect 8430 28906 8580 28920
rect 8430 27734 8460 28906
rect 8700 28906 8850 28920
rect 8820 28334 8850 28906
rect 8700 28320 8850 28334
rect 8910 28906 9090 28920
rect 8910 28334 8940 28906
rect 9060 28334 9090 28906
rect 8910 28320 9090 28334
rect 9150 28906 9300 28920
rect 9150 28334 9180 28906
rect 9150 28320 9300 28334
rect 9420 28906 9570 28920
rect 8430 27720 8580 27734
rect 9540 27734 9570 28906
rect 9420 27720 9570 27734
rect 9630 28860 9840 28920
rect 9630 27990 9674 28860
rect 9796 27990 9840 28860
rect 9630 27720 9840 27990
rect 9900 27720 9990 28920
rect 10050 28906 10350 28920
rect 10050 27734 10140 28906
rect 10260 27734 10350 28906
rect 10050 27720 10350 27734
rect 10410 27720 10500 28920
rect 10560 28860 10770 28920
rect 10560 27990 10604 28860
rect 10726 27990 10770 28860
rect 10560 27720 10770 27990
rect 10830 28906 10980 28920
rect 10830 27734 10860 28906
rect 10830 27720 10980 27734
rect 11100 28906 11250 28920
rect 11220 27734 11250 28906
rect 11100 27720 11250 27734
rect 11310 27720 11400 28920
rect 11460 28906 11640 28920
rect 11460 27734 11490 28906
rect 11610 28320 11640 28906
rect 11700 28906 11850 28920
rect 11700 28334 11730 28906
rect 11700 28320 11850 28334
rect 12060 28906 12210 28920
rect 12180 28334 12210 28906
rect 12060 28320 12210 28334
rect 12270 28906 12450 28920
rect 12270 28334 12300 28906
rect 12420 28334 12450 28906
rect 12270 28320 12450 28334
rect 12510 28906 12660 28920
rect 12510 28334 12540 28906
rect 12510 28320 12660 28334
rect 12780 28906 12930 28920
rect 12900 28334 12930 28906
rect 12780 28320 12930 28334
rect 12990 28906 13170 28920
rect 12990 28334 13020 28906
rect 13140 28334 13170 28906
rect 12990 28320 13170 28334
rect 13230 28906 13380 28920
rect 13230 28334 13260 28906
rect 13230 28320 13380 28334
rect 13740 28906 13890 28920
rect 13860 28334 13890 28906
rect 13740 28320 13890 28334
rect 13950 28906 14130 28920
rect 13950 28334 13980 28906
rect 14100 28334 14130 28906
rect 13950 28320 14130 28334
rect 14190 28906 14370 28920
rect 14190 28334 14220 28906
rect 14340 28334 14370 28906
rect 14190 28320 14370 28334
rect 14430 28906 14580 28920
rect 14430 28334 14460 28906
rect 14430 28320 14580 28334
rect 15420 28906 15570 28920
rect 15540 28334 15570 28906
rect 15420 28320 15570 28334
rect 15630 28906 15810 28920
rect 15630 28334 15660 28906
rect 15780 28334 15810 28906
rect 15630 28320 15810 28334
rect 15870 28906 16020 28920
rect 15870 28334 15900 28906
rect 15870 28320 16020 28334
rect 16620 28906 16770 28920
rect 16740 28334 16770 28906
rect 16620 28320 16770 28334
rect 16830 28906 17010 28920
rect 16830 28334 16860 28906
rect 16980 28334 17010 28906
rect 16830 28320 17010 28334
rect 17070 28906 17220 28920
rect 17070 28334 17100 28906
rect 17070 28320 17220 28334
rect 18060 28906 18210 28920
rect 18180 28334 18210 28906
rect 18060 28320 18210 28334
rect 18270 28906 18450 28920
rect 18270 28334 18300 28906
rect 18420 28334 18450 28906
rect 18270 28320 18450 28334
rect 18510 28906 18660 28920
rect 18510 28334 18540 28906
rect 18510 28320 18660 28334
rect 19350 28906 19500 28920
rect 19470 28334 19500 28906
rect 19350 28320 19500 28334
rect 19560 28906 19740 28920
rect 19560 28320 19590 28906
rect 11460 27720 11610 27734
rect 19710 27734 19740 28906
rect 19590 27720 19740 27734
rect 19800 27720 19890 28920
rect 19950 28906 20100 28920
rect 19950 27734 19980 28906
rect 20940 28906 21090 28920
rect 21060 28334 21090 28906
rect 20940 28320 21090 28334
rect 21150 28906 21330 28920
rect 21150 28334 21180 28906
rect 21300 28334 21330 28906
rect 21150 28320 21330 28334
rect 21390 28906 21540 28920
rect 21390 28334 21420 28906
rect 21390 28320 21540 28334
rect 22140 28906 22290 28920
rect 22260 28334 22290 28906
rect 22140 28320 22290 28334
rect 22350 28906 22530 28920
rect 22350 28334 22380 28906
rect 22500 28334 22530 28906
rect 22350 28320 22530 28334
rect 22590 28906 22740 28920
rect 22590 28334 22620 28906
rect 22590 28320 22740 28334
rect 23580 28906 23730 28920
rect 23700 28334 23730 28906
rect 23580 28320 23730 28334
rect 23790 28906 23970 28920
rect 23790 28334 23820 28906
rect 23940 28334 23970 28906
rect 23790 28320 23970 28334
rect 24030 28906 24180 28920
rect 24030 28334 24060 28906
rect 24030 28320 24180 28334
rect 25020 28906 25170 28920
rect 25140 28334 25170 28906
rect 25020 28320 25170 28334
rect 25230 28906 25410 28920
rect 25230 28334 25260 28906
rect 25380 28334 25410 28906
rect 25230 28320 25410 28334
rect 25470 28906 25620 28920
rect 25470 28334 25500 28906
rect 25470 28320 25620 28334
rect 26460 28906 26610 28920
rect 26580 28334 26610 28906
rect 26460 28320 26610 28334
rect 26670 28906 26850 28920
rect 26670 28334 26700 28906
rect 26820 28334 26850 28906
rect 26670 28320 26850 28334
rect 26910 28906 27060 28920
rect 26910 28334 26940 28906
rect 26910 28320 27060 28334
rect 28470 28906 28620 28920
rect 28590 28334 28620 28906
rect 28470 28320 28620 28334
rect 28680 28906 28860 28920
rect 28680 28320 28710 28906
rect 19950 27720 20100 27734
rect 28830 27734 28860 28906
rect 28710 27720 28860 27734
rect 28920 27720 29010 28920
rect 29070 28906 29220 28920
rect 29070 27734 29100 28906
rect 30300 28906 30450 28920
rect 30420 28334 30450 28906
rect 30300 28320 30450 28334
rect 30510 28906 30690 28920
rect 30510 28334 30540 28906
rect 30660 28334 30690 28906
rect 30510 28320 30690 28334
rect 30750 28906 30900 28920
rect 30750 28334 30780 28906
rect 30750 28320 30900 28334
rect 31830 28906 31980 28920
rect 31950 28334 31980 28906
rect 31830 28320 31980 28334
rect 32040 28906 32220 28920
rect 32040 28320 32070 28906
rect 29070 27720 29220 27734
rect 32190 27734 32220 28906
rect 32070 27720 32220 27734
rect 32280 27720 32370 28920
rect 32430 28906 32580 28920
rect 32430 27734 32460 28906
rect 32430 27720 32580 27734
rect 32940 28906 33090 28920
rect 33060 27734 33090 28906
rect 32940 27720 33090 27734
rect 33150 28860 33360 28920
rect 33150 27990 33194 28860
rect 33316 27990 33360 28860
rect 33150 27720 33360 27990
rect 33420 27720 33510 28920
rect 33570 28906 33870 28920
rect 33570 27734 33660 28906
rect 33780 27734 33870 28906
rect 33570 27720 33870 27734
rect 33930 27720 34020 28920
rect 34080 28860 34290 28920
rect 34080 27990 34124 28860
rect 34246 27990 34290 28860
rect 34080 27720 34290 27990
rect 34350 28906 34500 28920
rect 34350 27734 34380 28906
rect 34860 28906 35010 28920
rect 34980 28334 35010 28906
rect 34860 28320 35010 28334
rect 35070 28906 35250 28920
rect 35070 28334 35100 28906
rect 35220 28334 35250 28906
rect 35070 28320 35250 28334
rect 35310 28906 35460 28920
rect 35310 28334 35340 28906
rect 35310 28320 35460 28334
rect 36060 28906 36210 28920
rect 36180 28334 36210 28906
rect 36060 28320 36210 28334
rect 36270 28906 36450 28920
rect 36270 28334 36300 28906
rect 36420 28334 36450 28906
rect 36270 28320 36450 28334
rect 36510 28906 36660 28920
rect 36510 28334 36540 28906
rect 36510 28320 36660 28334
rect 37500 28906 37650 28920
rect 37620 28334 37650 28906
rect 37500 28320 37650 28334
rect 37710 28906 37890 28920
rect 37710 28334 37740 28906
rect 37860 28334 37890 28906
rect 37710 28320 37890 28334
rect 37950 28906 38100 28920
rect 37950 28334 37980 28906
rect 37950 28320 38100 28334
rect 38700 28906 38850 28920
rect 38820 28334 38850 28906
rect 38700 28320 38850 28334
rect 38910 28906 39090 28920
rect 38910 28334 38940 28906
rect 39060 28334 39090 28906
rect 38910 28320 39090 28334
rect 39150 28906 39300 28920
rect 39150 28334 39180 28906
rect 39150 28320 39300 28334
rect 39660 28906 39810 28920
rect 34350 27720 34500 27734
rect 39780 27734 39810 28906
rect 39660 27720 39810 27734
rect 39870 28860 40080 28920
rect 39870 27990 39914 28860
rect 40036 27990 40080 28860
rect 39870 27720 40080 27990
rect 40140 27720 40230 28920
rect 40290 28906 40590 28920
rect 40290 27734 40380 28906
rect 40500 27734 40590 28906
rect 40290 27720 40590 27734
rect 40650 27720 40740 28920
rect 40800 28860 41010 28920
rect 40800 27990 40844 28860
rect 40966 27990 41010 28860
rect 40800 27720 41010 27990
rect 41070 28906 41220 28920
rect 41070 27734 41100 28906
rect 41580 28906 41730 28920
rect 41700 28334 41730 28906
rect 41580 28320 41730 28334
rect 41790 28906 41970 28920
rect 41790 28334 41820 28906
rect 41940 28334 41970 28906
rect 41790 28320 41970 28334
rect 42030 28906 42180 28920
rect 42030 28334 42060 28906
rect 42030 28320 42180 28334
rect 43110 28906 43260 28920
rect 43230 28334 43260 28906
rect 43110 28320 43260 28334
rect 43320 28906 43500 28920
rect 43320 28320 43350 28906
rect 41070 27720 41220 27734
rect 43470 27734 43500 28906
rect 43350 27720 43500 27734
rect 43560 27720 43650 28920
rect 43710 28906 43860 28920
rect 43710 27734 43740 28906
rect 43710 27720 43860 27734
rect 44460 28906 44610 28920
rect 44580 27734 44610 28906
rect 44460 27720 44610 27734
rect 44670 27720 44760 28920
rect 44820 28906 45000 28920
rect 44820 27734 44850 28906
rect 44970 28320 45000 28906
rect 45060 28906 45210 28920
rect 45060 28334 45090 28906
rect 45060 28320 45210 28334
rect 45900 28906 46050 28920
rect 44820 27720 44970 27734
rect 46020 27734 46050 28906
rect 45900 27720 46050 27734
rect 46110 27720 46200 28920
rect 46260 28906 46440 28920
rect 46260 27734 46290 28906
rect 46410 28320 46440 28906
rect 46500 28906 46650 28920
rect 46500 28334 46530 28906
rect 46500 28320 46650 28334
rect 46860 28890 47010 28920
rect 46980 28320 47010 28890
rect 47070 28890 47220 28920
rect 47070 28320 47100 28890
rect 47340 28906 47490 28920
rect 46260 27720 46410 27734
rect 47460 27734 47490 28906
rect 47340 27720 47490 27734
rect 47550 28740 47730 28920
rect 47550 27720 47580 28740
rect 47700 27720 47730 28740
rect 47790 28906 47970 28920
rect 47790 27734 47820 28906
rect 47940 27734 47970 28906
rect 47790 27720 47970 27734
rect 48030 27900 48060 28920
rect 48180 27900 48210 28920
rect 48030 27720 48210 27900
rect 48270 28876 48420 28920
rect 48270 27854 48300 28876
rect 48540 28906 48690 28920
rect 48660 28334 48690 28906
rect 48540 28320 48690 28334
rect 48750 28906 48930 28920
rect 48750 28334 48780 28906
rect 48900 28334 48930 28906
rect 48750 28320 48930 28334
rect 48990 28906 49140 28920
rect 48990 28334 49020 28906
rect 48990 28320 49140 28334
rect 49260 28906 49410 28920
rect 48270 27720 48420 27854
rect 49380 27734 49410 28906
rect 49260 27720 49410 27734
rect 49470 27720 49560 28920
rect 49620 28906 49800 28920
rect 49620 27734 49650 28906
rect 49770 28320 49800 28906
rect 49860 28906 50010 28920
rect 49860 28334 49890 28906
rect 49860 28320 50010 28334
rect 49620 27720 49770 27734
rect 5340 24466 5490 24480
rect 5460 23294 5490 24466
rect 5340 23280 5490 23294
rect 5550 24210 5760 24480
rect 5550 23340 5594 24210
rect 5716 23340 5760 24210
rect 5550 23280 5760 23340
rect 5820 23280 5910 24480
rect 5970 24466 6270 24480
rect 5970 23294 6060 24466
rect 6180 23294 6270 24466
rect 5970 23280 6270 23294
rect 6330 23280 6420 24480
rect 6480 24210 6690 24480
rect 6480 23340 6524 24210
rect 6646 23340 6690 24210
rect 6480 23280 6690 23340
rect 6750 24466 6900 24480
rect 6750 23294 6780 24466
rect 8070 24466 8220 24480
rect 6750 23280 6900 23294
rect 7020 23866 7170 23880
rect 7140 23294 7170 23866
rect 7020 23280 7170 23294
rect 7230 23866 7410 23880
rect 7230 23294 7260 23866
rect 7380 23294 7410 23866
rect 7230 23280 7410 23294
rect 7470 23866 7620 23880
rect 7470 23294 7500 23866
rect 7470 23280 7620 23294
rect 7830 23866 7980 23880
rect 7950 23294 7980 23866
rect 7830 23280 7980 23294
rect 8040 23294 8070 23880
rect 8190 23294 8220 24466
rect 8040 23280 8220 23294
rect 8280 23280 8370 24480
rect 8430 24466 8580 24480
rect 8430 23294 8460 24466
rect 9420 24466 9570 24480
rect 8430 23280 8580 23294
rect 8700 23866 8850 23880
rect 8820 23294 8850 23866
rect 8700 23280 8850 23294
rect 8910 23866 9090 23880
rect 8910 23294 8940 23866
rect 9060 23294 9090 23866
rect 8910 23280 9090 23294
rect 9150 23866 9300 23880
rect 9150 23294 9180 23866
rect 9150 23280 9300 23294
rect 9540 23294 9570 24466
rect 9420 23280 9570 23294
rect 9630 24210 9840 24480
rect 9630 23340 9674 24210
rect 9796 23340 9840 24210
rect 9630 23280 9840 23340
rect 9900 23280 9990 24480
rect 10050 24466 10350 24480
rect 10050 23294 10140 24466
rect 10260 23294 10350 24466
rect 10050 23280 10350 23294
rect 10410 23280 10500 24480
rect 10560 24210 10770 24480
rect 10560 23340 10604 24210
rect 10726 23340 10770 24210
rect 10560 23280 10770 23340
rect 10830 24466 10980 24480
rect 10830 23294 10860 24466
rect 10830 23280 10980 23294
rect 12060 24466 12210 24480
rect 12180 23294 12210 24466
rect 12060 23280 12210 23294
rect 12270 24466 12450 24480
rect 12270 23294 12300 24466
rect 12420 23294 12450 24466
rect 12270 23280 12450 23294
rect 12510 24300 12690 24480
rect 12510 23280 12540 24300
rect 12660 23280 12690 24300
rect 12750 24346 12900 24480
rect 12750 23324 12780 24346
rect 15270 24466 15420 24480
rect 12750 23280 12900 23324
rect 13860 23310 13890 23880
rect 13740 23280 13890 23310
rect 13950 23310 13980 23880
rect 13950 23280 14100 23310
rect 15030 23866 15180 23880
rect 15150 23294 15180 23866
rect 15030 23280 15180 23294
rect 15240 23294 15270 23880
rect 15390 23294 15420 24466
rect 15240 23280 15420 23294
rect 15480 23280 15570 24480
rect 15630 24466 15780 24480
rect 15630 23294 15660 24466
rect 25500 24466 25650 24480
rect 15630 23280 15780 23294
rect 20700 23866 20850 23880
rect 20820 23294 20850 23866
rect 20700 23280 20850 23294
rect 20910 23866 21090 23880
rect 20910 23294 20940 23866
rect 21060 23294 21090 23866
rect 20910 23280 21090 23294
rect 21150 23866 21300 23880
rect 21150 23294 21180 23866
rect 21150 23280 21300 23294
rect 23100 23866 23250 23880
rect 23220 23294 23250 23866
rect 23100 23280 23250 23294
rect 23310 23866 23490 23880
rect 23310 23294 23340 23866
rect 23460 23294 23490 23866
rect 23310 23280 23490 23294
rect 23550 23866 23700 23880
rect 23550 23294 23580 23866
rect 23550 23280 23700 23294
rect 25620 23294 25650 24466
rect 25500 23280 25650 23294
rect 25710 24210 25920 24480
rect 25710 23340 25754 24210
rect 25876 23340 25920 24210
rect 25710 23280 25920 23340
rect 25980 23280 26070 24480
rect 26130 24466 26430 24480
rect 26130 23294 26220 24466
rect 26340 23294 26430 24466
rect 26130 23280 26430 23294
rect 26490 23280 26580 24480
rect 26640 24210 26850 24480
rect 26640 23340 26684 24210
rect 26806 23340 26850 24210
rect 26640 23280 26850 23340
rect 26910 24466 27060 24480
rect 26910 23294 26940 24466
rect 28230 24466 28380 24480
rect 26910 23280 27060 23294
rect 27990 23866 28140 23880
rect 28110 23294 28140 23866
rect 27990 23280 28140 23294
rect 28200 23294 28230 23880
rect 28350 23294 28380 24466
rect 28200 23280 28380 23294
rect 28440 23280 28530 24480
rect 28590 24466 28740 24480
rect 28590 23294 28620 24466
rect 31350 24466 31500 24480
rect 28590 23280 28740 23294
rect 30420 23310 30450 23880
rect 30300 23280 30450 23310
rect 30510 23310 30540 23880
rect 30510 23280 30660 23310
rect 31110 23866 31260 23880
rect 31230 23294 31260 23866
rect 31110 23280 31260 23294
rect 31320 23294 31350 23880
rect 31470 23294 31500 24466
rect 31320 23280 31500 23294
rect 31560 23280 31650 24480
rect 31710 24466 31860 24480
rect 31710 23294 31740 24466
rect 31710 23280 31860 23294
rect 32340 23310 32370 23880
rect 32220 23280 32370 23310
rect 32430 23310 32460 23880
rect 32430 23280 32580 23310
rect 33180 23866 33330 23880
rect 33300 23294 33330 23866
rect 33180 23280 33330 23294
rect 33390 23866 33570 23880
rect 33390 23294 33420 23866
rect 33540 23294 33570 23866
rect 33390 23280 33570 23294
rect 33630 23866 33780 23880
rect 33630 23294 33660 23866
rect 33630 23280 33780 23294
rect 34620 23866 34770 23880
rect 34740 23294 34770 23866
rect 34620 23280 34770 23294
rect 34830 23866 35010 23880
rect 34830 23294 34860 23866
rect 34980 23294 35010 23866
rect 34830 23280 35010 23294
rect 35070 23866 35220 23880
rect 35070 23294 35100 23866
rect 35070 23280 35220 23294
rect 36060 23866 36210 23880
rect 36180 23294 36210 23866
rect 36060 23280 36210 23294
rect 36270 23866 36450 23880
rect 36270 23294 36300 23866
rect 36420 23294 36450 23866
rect 36270 23280 36450 23294
rect 36510 23866 36660 23880
rect 36510 23294 36540 23866
rect 36510 23280 36660 23294
rect 37500 23866 37650 23880
rect 37620 23294 37650 23866
rect 37500 23280 37650 23294
rect 37710 23866 37890 23880
rect 37710 23294 37740 23866
rect 37860 23294 37890 23866
rect 37710 23280 37890 23294
rect 37950 23866 38100 23880
rect 37950 23294 37980 23866
rect 37950 23280 38100 23294
rect 38940 23866 39090 23880
rect 39060 23294 39090 23866
rect 38940 23280 39090 23294
rect 39150 23866 39330 23880
rect 39150 23294 39180 23866
rect 39300 23294 39330 23866
rect 39150 23280 39330 23294
rect 39390 23866 39540 23880
rect 39390 23294 39420 23866
rect 39390 23280 39540 23294
rect 40380 23866 40530 23880
rect 40500 23294 40530 23866
rect 40380 23280 40530 23294
rect 40590 23866 40770 23880
rect 40590 23294 40620 23866
rect 40740 23294 40770 23866
rect 40590 23280 40770 23294
rect 40830 23866 40980 23880
rect 40830 23294 40860 23866
rect 40830 23280 40980 23294
rect 41820 23866 41970 23880
rect 41940 23294 41970 23866
rect 41820 23280 41970 23294
rect 42030 23866 42210 23880
rect 42030 23294 42060 23866
rect 42180 23294 42210 23866
rect 42030 23280 42210 23294
rect 42270 23866 42420 23880
rect 42270 23294 42300 23866
rect 42270 23280 42420 23294
rect 43380 23310 43410 24480
rect 43260 23280 43410 23310
rect 43470 23280 43560 24480
rect 43620 23310 43650 24480
rect 47820 24466 47970 24480
rect 43620 23280 43770 23310
rect 44580 23310 44610 23880
rect 44460 23280 44610 23310
rect 44670 23310 44700 23880
rect 44670 23280 44820 23310
rect 47940 23294 47970 24466
rect 47820 23280 47970 23294
rect 48030 24210 48240 24480
rect 48030 23340 48074 24210
rect 48196 23340 48240 24210
rect 48030 23280 48240 23340
rect 48300 23280 48390 24480
rect 48450 24466 48750 24480
rect 48450 23294 48540 24466
rect 48660 23294 48750 24466
rect 48450 23280 48750 23294
rect 48810 23280 48900 24480
rect 48960 24210 49170 24480
rect 48960 23340 49004 24210
rect 49126 23340 49170 24210
rect 48960 23280 49170 23340
rect 49230 24466 49380 24480
rect 49230 23294 49260 24466
rect 49230 23280 49380 23294
rect 5340 22906 5490 22920
rect 5460 21734 5490 22906
rect 5340 21720 5490 21734
rect 5550 22860 5760 22920
rect 5550 21990 5594 22860
rect 5716 21990 5760 22860
rect 5550 21720 5760 21990
rect 5820 21720 5910 22920
rect 5970 22906 6270 22920
rect 5970 21734 6060 22906
rect 6180 21734 6270 22906
rect 5970 21720 6270 21734
rect 6330 21720 6420 22920
rect 6480 22860 6690 22920
rect 6480 21990 6524 22860
rect 6646 21990 6690 22860
rect 6480 21720 6690 21990
rect 6750 22906 6900 22920
rect 6750 21734 6780 22906
rect 8220 22906 8370 22920
rect 8340 22334 8370 22906
rect 8220 22320 8370 22334
rect 8430 22906 8610 22920
rect 8430 22334 8460 22906
rect 8580 22334 8610 22906
rect 8430 22320 8610 22334
rect 8670 22906 8820 22920
rect 8670 22334 8700 22906
rect 8670 22320 8820 22334
rect 9660 22906 9810 22920
rect 9780 22334 9810 22906
rect 9660 22320 9810 22334
rect 9870 22906 10050 22920
rect 9870 22334 9900 22906
rect 10020 22334 10050 22906
rect 9870 22320 10050 22334
rect 10110 22906 10260 22920
rect 10110 22334 10140 22906
rect 10110 22320 10260 22334
rect 11190 22906 11340 22920
rect 11310 22334 11340 22906
rect 11190 22320 11340 22334
rect 11400 22906 11580 22920
rect 11400 22320 11430 22906
rect 6750 21720 6900 21734
rect 11550 21734 11580 22906
rect 11430 21720 11580 21734
rect 11640 21720 11730 22920
rect 11790 22906 11940 22920
rect 11790 21734 11820 22906
rect 11790 21720 11940 21734
rect 14220 22906 14370 22920
rect 14340 21734 14370 22906
rect 14220 21720 14370 21734
rect 14430 22860 14640 22920
rect 14430 21990 14474 22860
rect 14596 21990 14640 22860
rect 14430 21720 14640 21990
rect 14700 21720 14790 22920
rect 14850 22906 15150 22920
rect 14850 21734 14940 22906
rect 15060 21734 15150 22906
rect 14850 21720 15150 21734
rect 15210 21720 15300 22920
rect 15360 22860 15570 22920
rect 15360 21990 15404 22860
rect 15526 21990 15570 22860
rect 15360 21720 15570 21990
rect 15630 22906 15780 22920
rect 15630 21734 15660 22906
rect 16860 22890 17010 22920
rect 16980 22320 17010 22890
rect 17070 22890 17220 22920
rect 17070 22320 17100 22890
rect 18060 22906 18210 22920
rect 18180 22334 18210 22906
rect 18060 22320 18210 22334
rect 18270 22906 18450 22920
rect 18270 22334 18300 22906
rect 18420 22334 18450 22906
rect 18270 22320 18450 22334
rect 18510 22906 18660 22920
rect 18510 22334 18540 22906
rect 18510 22320 18660 22334
rect 18780 22906 18930 22920
rect 15630 21720 15780 21734
rect 18900 21734 18930 22906
rect 18780 21720 18930 21734
rect 18990 22860 19200 22920
rect 18990 21990 19034 22860
rect 19156 21990 19200 22860
rect 18990 21720 19200 21990
rect 19260 21720 19350 22920
rect 19410 22906 19710 22920
rect 19410 21734 19500 22906
rect 19620 21734 19710 22906
rect 19410 21720 19710 21734
rect 19770 21720 19860 22920
rect 19920 22860 20130 22920
rect 19920 21990 19964 22860
rect 20086 21990 20130 22860
rect 19920 21720 20130 21990
rect 20190 22906 20340 22920
rect 20190 21734 20220 22906
rect 20190 21720 20340 21734
rect 20460 22906 20610 22920
rect 20580 21734 20610 22906
rect 20460 21720 20610 21734
rect 20670 22860 20880 22920
rect 20670 21990 20714 22860
rect 20836 21990 20880 22860
rect 20670 21720 20880 21990
rect 20940 21720 21030 22920
rect 21090 22906 21390 22920
rect 21090 21734 21180 22906
rect 21300 21734 21390 22906
rect 21090 21720 21390 21734
rect 21450 21720 21540 22920
rect 21600 22860 21810 22920
rect 21600 21990 21644 22860
rect 21766 21990 21810 22860
rect 21600 21720 21810 21990
rect 21870 22906 22020 22920
rect 21870 21734 21900 22906
rect 22230 22906 22380 22920
rect 22350 22334 22380 22906
rect 22230 22320 22380 22334
rect 22440 22906 22620 22920
rect 22440 22320 22470 22906
rect 21870 21720 22020 21734
rect 22590 21734 22620 22906
rect 22470 21720 22620 21734
rect 22680 21720 22770 22920
rect 22830 22906 22980 22920
rect 22830 21734 22860 22906
rect 25020 22890 25170 22920
rect 25140 22320 25170 22890
rect 25230 22890 25380 22920
rect 25230 22320 25260 22890
rect 26310 22906 26460 22920
rect 26430 22334 26460 22906
rect 26310 22320 26460 22334
rect 26520 22906 26700 22920
rect 26520 22320 26550 22906
rect 22830 21720 22980 21734
rect 26670 21734 26700 22906
rect 26550 21720 26700 21734
rect 26760 21720 26850 22920
rect 26910 22906 27060 22920
rect 26910 21734 26940 22906
rect 27990 22906 28140 22920
rect 28110 22334 28140 22906
rect 27990 22320 28140 22334
rect 28200 22906 28380 22920
rect 28200 22320 28230 22906
rect 26910 21720 27060 21734
rect 28350 21734 28380 22906
rect 28230 21720 28380 21734
rect 28440 21720 28530 22920
rect 28590 22906 28740 22920
rect 28590 21734 28620 22906
rect 29100 22906 29250 22920
rect 29220 22334 29250 22906
rect 29100 22320 29250 22334
rect 29310 22906 29490 22920
rect 29310 22334 29340 22906
rect 29460 22334 29490 22906
rect 29310 22320 29490 22334
rect 29550 22906 29700 22920
rect 29550 22334 29580 22906
rect 29550 22320 29700 22334
rect 30300 22906 30450 22920
rect 28590 21720 28740 21734
rect 30420 21734 30450 22906
rect 30300 21720 30450 21734
rect 30510 21720 30600 22920
rect 30660 22906 30840 22920
rect 30660 21734 30690 22906
rect 30810 22320 30840 22906
rect 30900 22906 31050 22920
rect 30900 22334 30930 22906
rect 30900 22320 31050 22334
rect 31980 22906 32130 22920
rect 32100 22334 32130 22906
rect 31980 22320 32130 22334
rect 32190 22906 32370 22920
rect 32190 22334 32220 22906
rect 32340 22334 32370 22906
rect 32190 22320 32370 22334
rect 32430 22906 32580 22920
rect 32430 22334 32460 22906
rect 32430 22320 32580 22334
rect 33180 22906 33330 22920
rect 33300 22334 33330 22906
rect 33180 22320 33330 22334
rect 33390 22906 33570 22920
rect 33390 22334 33420 22906
rect 33540 22334 33570 22906
rect 33390 22320 33570 22334
rect 33630 22906 33780 22920
rect 33630 22334 33660 22906
rect 33630 22320 33780 22334
rect 34620 22906 34770 22920
rect 34740 22334 34770 22906
rect 34620 22320 34770 22334
rect 34830 22906 35010 22920
rect 34830 22334 34860 22906
rect 34980 22334 35010 22906
rect 34830 22320 35010 22334
rect 35070 22906 35220 22920
rect 35070 22334 35100 22906
rect 35070 22320 35220 22334
rect 35820 22906 35970 22920
rect 35940 22334 35970 22906
rect 35820 22320 35970 22334
rect 36030 22906 36210 22920
rect 36030 22334 36060 22906
rect 36180 22334 36210 22906
rect 36030 22320 36210 22334
rect 36270 22906 36420 22920
rect 36270 22334 36300 22906
rect 36270 22320 36420 22334
rect 36780 22906 36930 22920
rect 30660 21720 30810 21734
rect 36900 21734 36930 22906
rect 36780 21720 36930 21734
rect 36990 22860 37200 22920
rect 36990 21990 37034 22860
rect 37156 21990 37200 22860
rect 36990 21720 37200 21990
rect 37260 21720 37350 22920
rect 37410 22906 37710 22920
rect 37410 21734 37500 22906
rect 37620 21734 37710 22906
rect 37410 21720 37710 21734
rect 37770 21720 37860 22920
rect 37920 22860 38130 22920
rect 37920 21990 37964 22860
rect 38086 21990 38130 22860
rect 37920 21720 38130 21990
rect 38190 22906 38340 22920
rect 38190 21734 38220 22906
rect 39030 22906 39180 22920
rect 39150 22334 39180 22906
rect 39030 22320 39180 22334
rect 39240 22906 39420 22920
rect 39240 22320 39270 22906
rect 38190 21720 38340 21734
rect 39390 21734 39420 22906
rect 39270 21720 39420 21734
rect 39480 21720 39570 22920
rect 39630 22906 39780 22920
rect 39630 21734 39660 22906
rect 40380 22906 40530 22920
rect 40500 22334 40530 22906
rect 40380 22320 40530 22334
rect 40590 22906 40770 22920
rect 40590 22334 40620 22906
rect 40740 22334 40770 22906
rect 40590 22320 40770 22334
rect 40830 22906 40980 22920
rect 40830 22334 40860 22906
rect 40830 22320 40980 22334
rect 41670 22906 41820 22920
rect 41790 22334 41820 22906
rect 41670 22320 41820 22334
rect 41880 22906 42060 22920
rect 41880 22320 41910 22906
rect 39630 21720 39780 21734
rect 42030 21734 42060 22906
rect 41910 21720 42060 21734
rect 42120 21720 42210 22920
rect 42270 22906 42420 22920
rect 42270 21734 42300 22906
rect 42270 21720 42420 21734
rect 43260 22890 43410 22920
rect 43380 21720 43410 22890
rect 43470 21720 43560 22920
rect 43620 22890 43770 22920
rect 43620 21720 43650 22890
rect 44220 22906 44370 22920
rect 44340 21734 44370 22906
rect 44220 21720 44370 21734
rect 44430 22860 44640 22920
rect 44430 21990 44474 22860
rect 44596 21990 44640 22860
rect 44430 21720 44640 21990
rect 44700 21720 44790 22920
rect 44850 22906 45150 22920
rect 44850 21734 44940 22906
rect 45060 21734 45150 22906
rect 44850 21720 45150 21734
rect 45210 21720 45300 22920
rect 45360 22860 45570 22920
rect 45360 21990 45404 22860
rect 45526 21990 45570 22860
rect 45360 21720 45570 21990
rect 45630 22906 45780 22920
rect 45630 21734 45660 22906
rect 45630 21720 45780 21734
rect 45900 22906 46050 22920
rect 46020 21734 46050 22906
rect 45900 21720 46050 21734
rect 46110 22860 46320 22920
rect 46110 21990 46154 22860
rect 46276 21990 46320 22860
rect 46110 21720 46320 21990
rect 46380 21720 46470 22920
rect 46530 22906 46830 22920
rect 46530 21734 46620 22906
rect 46740 21734 46830 22906
rect 46530 21720 46830 21734
rect 46890 21720 46980 22920
rect 47040 22860 47250 22920
rect 47040 21990 47084 22860
rect 47206 21990 47250 22860
rect 47040 21720 47250 21990
rect 47310 22906 47460 22920
rect 47310 21734 47340 22906
rect 47580 22890 47730 22920
rect 47700 22320 47730 22890
rect 47790 22890 47940 22920
rect 47790 22320 47820 22890
rect 48780 22906 48930 22920
rect 47310 21720 47460 21734
rect 48900 21734 48930 22906
rect 48780 21720 48930 21734
rect 48990 22740 49170 22920
rect 48990 21720 49020 22740
rect 49140 21720 49170 22740
rect 49230 22906 49410 22920
rect 49230 21734 49260 22906
rect 49380 21734 49410 22906
rect 49230 21720 49410 21734
rect 49470 21900 49500 22920
rect 49620 21900 49650 22920
rect 49470 21720 49650 21900
rect 49710 22876 49860 22920
rect 49710 21854 49740 22876
rect 49710 21720 49860 21854
rect 5910 18466 6060 18480
rect 5670 17866 5820 17880
rect 5790 17294 5820 17866
rect 5670 17280 5820 17294
rect 5880 17294 5910 17880
rect 6030 17294 6060 18466
rect 5880 17280 6060 17294
rect 6120 17280 6210 18480
rect 6270 18466 6420 18480
rect 6270 17294 6300 18466
rect 6270 17280 6420 17294
rect 8940 18466 9090 18480
rect 9060 17294 9090 18466
rect 8940 17280 9090 17294
rect 9150 18210 9360 18480
rect 9150 17340 9194 18210
rect 9316 17340 9360 18210
rect 9150 17280 9360 17340
rect 9420 17280 9510 18480
rect 9570 18466 9870 18480
rect 9570 17294 9660 18466
rect 9780 17294 9870 18466
rect 9570 17280 9870 17294
rect 9930 17280 10020 18480
rect 10080 18210 10290 18480
rect 10080 17340 10124 18210
rect 10246 17340 10290 18210
rect 10080 17280 10290 17340
rect 10350 18466 10500 18480
rect 10350 17294 10380 18466
rect 10350 17280 10500 17294
rect 11580 18466 11730 18480
rect 11700 17294 11730 18466
rect 11580 17280 11730 17294
rect 11790 18210 12000 18480
rect 11790 17340 11834 18210
rect 11956 17340 12000 18210
rect 11790 17280 12000 17340
rect 12060 17280 12150 18480
rect 12210 18466 12510 18480
rect 12210 17294 12300 18466
rect 12420 17294 12510 18466
rect 12210 17280 12510 17294
rect 12570 17280 12660 18480
rect 12720 18210 12930 18480
rect 12720 17340 12764 18210
rect 12886 17340 12930 18210
rect 12720 17280 12930 17340
rect 12990 18466 13140 18480
rect 12990 17294 13020 18466
rect 12990 17280 13140 17294
rect 13500 18466 13650 18480
rect 13620 17294 13650 18466
rect 13500 17280 13650 17294
rect 13710 18210 13920 18480
rect 13710 17340 13754 18210
rect 13876 17340 13920 18210
rect 13710 17280 13920 17340
rect 13980 17280 14070 18480
rect 14130 18466 14430 18480
rect 14130 17294 14220 18466
rect 14340 17294 14430 18466
rect 14130 17280 14430 17294
rect 14490 17280 14580 18480
rect 14640 18210 14850 18480
rect 14640 17340 14684 18210
rect 14806 17340 14850 18210
rect 14640 17280 14850 17340
rect 14910 18466 15060 18480
rect 14910 17294 14940 18466
rect 14910 17280 15060 17294
rect 15420 18346 15570 18480
rect 15540 17324 15570 18346
rect 15420 17280 15570 17324
rect 15630 18300 15810 18480
rect 15630 17280 15660 18300
rect 15780 17280 15810 18300
rect 15870 18466 16050 18480
rect 15870 17294 15900 18466
rect 16020 17294 16050 18466
rect 15870 17280 16050 17294
rect 16110 18466 16260 18480
rect 16110 17294 16140 18466
rect 18150 18466 18300 18480
rect 16110 17280 16260 17294
rect 17910 17866 18060 17880
rect 18030 17294 18060 17866
rect 17910 17280 18060 17294
rect 18120 17294 18150 17880
rect 18270 17294 18300 18466
rect 18120 17280 18300 17294
rect 18360 17280 18450 18480
rect 18510 18466 18660 18480
rect 18510 17294 18540 18466
rect 24540 18466 24690 18480
rect 18510 17280 18660 17294
rect 19500 17866 19650 17880
rect 19620 17294 19650 17866
rect 19500 17280 19650 17294
rect 19710 17866 19890 17880
rect 19710 17294 19740 17866
rect 19860 17294 19890 17866
rect 19710 17280 19890 17294
rect 19950 17866 20100 17880
rect 19950 17294 19980 17866
rect 19950 17280 20100 17294
rect 20940 17866 21090 17880
rect 21060 17294 21090 17866
rect 20940 17280 21090 17294
rect 21150 17866 21330 17880
rect 21150 17294 21180 17866
rect 21300 17294 21330 17866
rect 21150 17280 21330 17294
rect 21390 17866 21540 17880
rect 21390 17294 21420 17866
rect 21390 17280 21540 17294
rect 22140 17866 22290 17880
rect 22260 17294 22290 17866
rect 22140 17280 22290 17294
rect 22350 17866 22530 17880
rect 22350 17294 22380 17866
rect 22500 17294 22530 17866
rect 22350 17280 22530 17294
rect 22590 17866 22740 17880
rect 22590 17294 22620 17866
rect 22590 17280 22740 17294
rect 23580 17866 23730 17880
rect 23700 17294 23730 17866
rect 23580 17280 23730 17294
rect 23790 17866 23970 17880
rect 23790 17294 23820 17866
rect 23940 17294 23970 17866
rect 23790 17280 23970 17294
rect 24030 17866 24180 17880
rect 24030 17294 24060 17866
rect 24030 17280 24180 17294
rect 24660 17294 24690 18466
rect 24540 17280 24690 17294
rect 24750 18210 24960 18480
rect 24750 17340 24794 18210
rect 24916 17340 24960 18210
rect 24750 17280 24960 17340
rect 25020 17280 25110 18480
rect 25170 18466 25470 18480
rect 25170 17294 25260 18466
rect 25380 17294 25470 18466
rect 25170 17280 25470 17294
rect 25530 17280 25620 18480
rect 25680 18210 25890 18480
rect 25680 17340 25724 18210
rect 25846 17340 25890 18210
rect 25680 17280 25890 17340
rect 25950 18466 26100 18480
rect 25950 17294 25980 18466
rect 25950 17280 26100 17294
rect 26220 18466 26370 18480
rect 26340 17294 26370 18466
rect 26220 17280 26370 17294
rect 26430 17280 26520 18480
rect 26580 18466 26730 18480
rect 26580 17294 26610 18466
rect 28710 18466 28860 18480
rect 26730 17294 26760 17880
rect 26580 17280 26760 17294
rect 26820 17866 26970 17880
rect 26820 17294 26850 17866
rect 26820 17280 26970 17294
rect 27300 17310 27330 17880
rect 27180 17280 27330 17310
rect 27390 17310 27420 17880
rect 27390 17280 27540 17310
rect 28470 17866 28620 17880
rect 28590 17294 28620 17866
rect 28470 17280 28620 17294
rect 28680 17294 28710 17880
rect 28830 17294 28860 18466
rect 28680 17280 28860 17294
rect 28920 17280 29010 18480
rect 29070 18466 29220 18480
rect 29070 17294 29100 18466
rect 33180 18466 33330 18480
rect 29070 17280 29220 17294
rect 30540 17866 30690 17880
rect 30660 17294 30690 17866
rect 30540 17280 30690 17294
rect 30750 17866 30930 17880
rect 30750 17294 30780 17866
rect 30900 17294 30930 17866
rect 30750 17280 30930 17294
rect 30990 17866 31140 17880
rect 30990 17294 31020 17866
rect 30990 17280 31140 17294
rect 31980 17866 32130 17880
rect 32100 17294 32130 17866
rect 31980 17280 32130 17294
rect 32190 17866 32370 17880
rect 32190 17294 32220 17866
rect 32340 17294 32370 17866
rect 32190 17280 32370 17294
rect 32430 17866 32580 17880
rect 32430 17294 32460 17866
rect 32430 17280 32580 17294
rect 33300 17294 33330 18466
rect 33180 17280 33330 17294
rect 33390 17280 33480 18480
rect 33540 18466 33690 18480
rect 33540 17294 33570 18466
rect 36780 18466 36930 18480
rect 33690 17294 33720 17880
rect 33540 17280 33720 17294
rect 33780 17866 33930 17880
rect 33780 17294 33810 17866
rect 33780 17280 33930 17294
rect 35820 17866 35970 17880
rect 35940 17294 35970 17866
rect 35820 17280 35970 17294
rect 36030 17866 36210 17880
rect 36030 17294 36060 17866
rect 36180 17294 36210 17866
rect 36030 17280 36210 17294
rect 36270 17866 36420 17880
rect 36270 17294 36300 17866
rect 36270 17280 36420 17294
rect 36900 17294 36930 18466
rect 36780 17280 36930 17294
rect 36990 18466 37170 18480
rect 36990 17294 37020 18466
rect 37140 17294 37170 18466
rect 36990 17280 37170 17294
rect 37230 18300 37410 18480
rect 37230 17280 37260 18300
rect 37380 17280 37410 18300
rect 37470 18346 37620 18480
rect 37470 17324 37500 18346
rect 42780 18346 42930 18480
rect 37470 17280 37620 17324
rect 37980 17866 38130 17880
rect 38100 17294 38130 17866
rect 37980 17280 38130 17294
rect 38190 17866 38370 17880
rect 38190 17294 38220 17866
rect 38340 17294 38370 17866
rect 38190 17280 38370 17294
rect 38430 17866 38580 17880
rect 38430 17294 38460 17866
rect 38430 17280 38580 17294
rect 38940 17866 39090 17880
rect 39060 17294 39090 17866
rect 38940 17280 39090 17294
rect 39150 17866 39330 17880
rect 39150 17294 39180 17866
rect 39300 17294 39330 17866
rect 39150 17280 39330 17294
rect 39390 17866 39540 17880
rect 39390 17294 39420 17866
rect 39390 17280 39540 17294
rect 40380 17866 40530 17880
rect 40500 17294 40530 17866
rect 40380 17280 40530 17294
rect 40590 17866 40770 17880
rect 40590 17294 40620 17866
rect 40740 17294 40770 17866
rect 40590 17280 40770 17294
rect 40830 17866 40980 17880
rect 40830 17294 40860 17866
rect 40830 17280 40980 17294
rect 41700 17310 41730 17880
rect 41580 17280 41730 17310
rect 41790 17310 41820 17880
rect 41790 17280 41940 17310
rect 42900 17324 42930 18346
rect 42780 17280 42930 17324
rect 42990 18300 43170 18480
rect 42990 17280 43020 18300
rect 43140 17280 43170 18300
rect 43230 18466 43410 18480
rect 43230 17294 43260 18466
rect 43380 17294 43410 18466
rect 43230 17280 43410 17294
rect 43470 17460 43500 18480
rect 43620 17460 43650 18480
rect 43470 17280 43650 17460
rect 43710 18466 43860 18480
rect 43710 17294 43740 18466
rect 43710 17280 43860 17294
rect 44460 18466 44610 18480
rect 44580 17294 44610 18466
rect 44460 17280 44610 17294
rect 44670 17280 44760 18480
rect 44820 18466 44970 18480
rect 44820 17294 44850 18466
rect 44970 17294 45000 17880
rect 44820 17280 45000 17294
rect 45060 17866 45210 17880
rect 45060 17294 45090 17866
rect 45060 17280 45210 17294
rect 46140 17866 46290 17880
rect 46260 17294 46290 17866
rect 46140 17280 46290 17294
rect 46350 17866 46530 17880
rect 46350 17294 46380 17866
rect 46500 17294 46530 17866
rect 46350 17280 46530 17294
rect 46590 17866 46740 17880
rect 46590 17294 46620 17866
rect 46590 17280 46740 17294
rect 47700 17310 47730 18480
rect 47580 17280 47730 17310
rect 47790 17280 47880 18480
rect 47940 17310 47970 18480
rect 47940 17280 48090 17310
rect 49020 18466 49170 18480
rect 49140 17294 49170 18466
rect 49020 17280 49170 17294
rect 49230 17280 49320 18480
rect 49380 18466 49530 18480
rect 49380 17294 49410 18466
rect 49530 17294 49560 17880
rect 49380 17280 49560 17294
rect 49620 17866 49770 17880
rect 49620 17294 49650 17866
rect 49620 17280 49770 17294
rect 6300 16906 6450 16920
rect 6420 16334 6450 16906
rect 6300 16320 6450 16334
rect 6510 16906 6690 16920
rect 6510 16334 6540 16906
rect 6660 16334 6690 16906
rect 6510 16320 6690 16334
rect 6750 16906 6900 16920
rect 6750 16334 6780 16906
rect 6750 16320 6900 16334
rect 7740 16906 7890 16920
rect 7860 15734 7890 16906
rect 7740 15720 7890 15734
rect 7950 16860 8160 16920
rect 7950 15990 7994 16860
rect 8116 15990 8160 16860
rect 7950 15720 8160 15990
rect 8220 15720 8310 16920
rect 8370 16906 8670 16920
rect 8370 15734 8460 16906
rect 8580 15734 8670 16906
rect 8370 15720 8670 15734
rect 8730 15720 8820 16920
rect 8880 16860 9090 16920
rect 8880 15990 8924 16860
rect 9046 15990 9090 16860
rect 8880 15720 9090 15990
rect 9150 16906 9300 16920
rect 9150 15734 9180 16906
rect 9150 15720 9300 15734
rect 9420 16906 9570 16920
rect 9540 15734 9570 16906
rect 9420 15720 9570 15734
rect 9630 16860 9840 16920
rect 9630 15990 9674 16860
rect 9796 15990 9840 16860
rect 9630 15720 9840 15990
rect 9900 15720 9990 16920
rect 10050 16906 10350 16920
rect 10050 15734 10140 16906
rect 10260 15734 10350 16906
rect 10050 15720 10350 15734
rect 10410 15720 10500 16920
rect 10560 16860 10770 16920
rect 10560 15990 10604 16860
rect 10726 15990 10770 16860
rect 10560 15720 10770 15990
rect 10830 16906 10980 16920
rect 10830 15734 10860 16906
rect 10830 15720 10980 15734
rect 11100 16906 11250 16920
rect 11220 15734 11250 16906
rect 11100 15720 11250 15734
rect 11310 16860 11520 16920
rect 11310 15990 11354 16860
rect 11476 15990 11520 16860
rect 11310 15720 11520 15990
rect 11580 15720 11670 16920
rect 11730 16906 12030 16920
rect 11730 15734 11820 16906
rect 11940 15734 12030 16906
rect 11730 15720 12030 15734
rect 12090 15720 12180 16920
rect 12240 16860 12450 16920
rect 12240 15990 12284 16860
rect 12406 15990 12450 16860
rect 12240 15720 12450 15990
rect 12510 16906 12660 16920
rect 12510 15734 12540 16906
rect 12510 15720 12660 15734
rect 13260 16906 13410 16920
rect 13380 15734 13410 16906
rect 13260 15720 13410 15734
rect 13470 16860 13680 16920
rect 13470 15990 13514 16860
rect 13636 15990 13680 16860
rect 13470 15720 13680 15990
rect 13740 15720 13830 16920
rect 13890 16906 14190 16920
rect 13890 15734 13980 16906
rect 14100 15734 14190 16906
rect 13890 15720 14190 15734
rect 14250 15720 14340 16920
rect 14400 16860 14610 16920
rect 14400 15990 14444 16860
rect 14566 15990 14610 16860
rect 14400 15720 14610 15990
rect 14670 16906 14820 16920
rect 14670 15734 14700 16906
rect 14670 15720 14820 15734
rect 14940 16906 15090 16920
rect 15060 15734 15090 16906
rect 14940 15720 15090 15734
rect 15150 16860 15360 16920
rect 15150 15990 15194 16860
rect 15316 15990 15360 16860
rect 15150 15720 15360 15990
rect 15420 15720 15510 16920
rect 15570 16906 15870 16920
rect 15570 15734 15660 16906
rect 15780 15734 15870 16906
rect 15570 15720 15870 15734
rect 15930 15720 16020 16920
rect 16080 16860 16290 16920
rect 16080 15990 16124 16860
rect 16246 15990 16290 16860
rect 16080 15720 16290 15990
rect 16350 16906 16500 16920
rect 16350 15734 16380 16906
rect 16350 15720 16500 15734
rect 16620 16876 16770 16920
rect 16740 15854 16770 16876
rect 16620 15720 16770 15854
rect 16830 15900 16860 16920
rect 16980 15900 17010 16920
rect 16830 15720 17010 15900
rect 17070 16906 17250 16920
rect 17070 15734 17100 16906
rect 17220 15734 17250 16906
rect 17070 15720 17250 15734
rect 17310 16906 17460 16920
rect 17310 15734 17340 16906
rect 17580 16890 17730 16920
rect 17700 16320 17730 16890
rect 17790 16890 17940 16920
rect 17790 16320 17820 16890
rect 18150 16906 18300 16920
rect 18270 16334 18300 16906
rect 18150 16320 18300 16334
rect 18360 16906 18540 16920
rect 18360 16320 18390 16906
rect 17310 15720 17460 15734
rect 18510 15734 18540 16906
rect 18390 15720 18540 15734
rect 18600 15720 18690 16920
rect 18750 16906 18900 16920
rect 18750 15734 18780 16906
rect 19260 16906 19410 16920
rect 19380 16334 19410 16906
rect 19260 16320 19410 16334
rect 19470 16906 19650 16920
rect 19470 16334 19500 16906
rect 19620 16334 19650 16906
rect 19470 16320 19650 16334
rect 19710 16906 19860 16920
rect 19710 16334 19740 16906
rect 19710 16320 19860 16334
rect 20700 16906 20850 16920
rect 18750 15720 18900 15734
rect 20820 15734 20850 16906
rect 20700 15720 20850 15734
rect 20910 15720 21000 16920
rect 21060 16906 21240 16920
rect 21060 15734 21090 16906
rect 21210 16320 21240 16906
rect 21300 16906 21450 16920
rect 21300 16334 21330 16906
rect 21300 16320 21450 16334
rect 22230 16906 22380 16920
rect 22350 16334 22380 16906
rect 22230 16320 22380 16334
rect 22440 16906 22620 16920
rect 22440 16320 22470 16906
rect 21060 15720 21210 15734
rect 22590 15734 22620 16906
rect 22470 15720 22620 15734
rect 22680 15720 22770 16920
rect 22830 16906 22980 16920
rect 22830 15734 22860 16906
rect 23580 16906 23730 16920
rect 23700 16334 23730 16906
rect 23580 16320 23730 16334
rect 23790 16906 23970 16920
rect 23790 16334 23820 16906
rect 23940 16334 23970 16906
rect 23790 16320 23970 16334
rect 24030 16906 24180 16920
rect 24030 16334 24060 16906
rect 24030 16320 24180 16334
rect 24780 16906 24930 16920
rect 24900 16334 24930 16906
rect 24780 16320 24930 16334
rect 24990 16906 25170 16920
rect 24990 16334 25020 16906
rect 25140 16334 25170 16906
rect 24990 16320 25170 16334
rect 25230 16906 25380 16920
rect 25230 16334 25260 16906
rect 25230 16320 25380 16334
rect 25740 16906 25890 16920
rect 22830 15720 22980 15734
rect 25860 15734 25890 16906
rect 25740 15720 25890 15734
rect 25950 16860 26160 16920
rect 25950 15990 25994 16860
rect 26116 15990 26160 16860
rect 25950 15720 26160 15990
rect 26220 15720 26310 16920
rect 26370 16906 26670 16920
rect 26370 15734 26460 16906
rect 26580 15734 26670 16906
rect 26370 15720 26670 15734
rect 26730 15720 26820 16920
rect 26880 16860 27090 16920
rect 26880 15990 26924 16860
rect 27046 15990 27090 16860
rect 26880 15720 27090 15990
rect 27150 16906 27300 16920
rect 27150 15734 27180 16906
rect 27900 16906 28050 16920
rect 28020 16334 28050 16906
rect 27900 16320 28050 16334
rect 28110 16906 28290 16920
rect 28110 16334 28140 16906
rect 28260 16334 28290 16906
rect 28110 16320 28290 16334
rect 28350 16906 28500 16920
rect 28350 16334 28380 16906
rect 28350 16320 28500 16334
rect 29100 16906 29250 16920
rect 29220 16334 29250 16906
rect 29100 16320 29250 16334
rect 29310 16906 29490 16920
rect 29310 16334 29340 16906
rect 29460 16334 29490 16906
rect 29310 16320 29490 16334
rect 29550 16906 29700 16920
rect 29550 16334 29580 16906
rect 29550 16320 29700 16334
rect 30300 16906 30450 16920
rect 27150 15720 27300 15734
rect 30420 15734 30450 16906
rect 30300 15720 30450 15734
rect 30510 16860 30720 16920
rect 30510 15990 30554 16860
rect 30676 15990 30720 16860
rect 30510 15720 30720 15990
rect 30780 15720 30870 16920
rect 30930 16906 31230 16920
rect 30930 15734 31020 16906
rect 31140 15734 31230 16906
rect 30930 15720 31230 15734
rect 31290 15720 31380 16920
rect 31440 16860 31650 16920
rect 31440 15990 31484 16860
rect 31606 15990 31650 16860
rect 31440 15720 31650 15990
rect 31710 16906 31860 16920
rect 31710 15734 31740 16906
rect 32220 16906 32370 16920
rect 32340 16334 32370 16906
rect 32220 16320 32370 16334
rect 32430 16906 32610 16920
rect 32430 16334 32460 16906
rect 32580 16334 32610 16906
rect 32430 16320 32610 16334
rect 32670 16906 32820 16920
rect 32670 16334 32700 16906
rect 32670 16320 32820 16334
rect 33180 16906 33330 16920
rect 33300 16334 33330 16906
rect 33180 16320 33330 16334
rect 33390 16906 33570 16920
rect 33390 16334 33420 16906
rect 33540 16334 33570 16906
rect 33390 16320 33570 16334
rect 33630 16906 33780 16920
rect 33630 16334 33660 16906
rect 33630 16320 33780 16334
rect 34620 16906 34770 16920
rect 34740 16334 34770 16906
rect 34620 16320 34770 16334
rect 34830 16906 35010 16920
rect 34830 16334 34860 16906
rect 34980 16334 35010 16906
rect 34830 16320 35010 16334
rect 35070 16906 35220 16920
rect 35070 16334 35100 16906
rect 35070 16320 35220 16334
rect 36060 16906 36210 16920
rect 31710 15720 31860 15734
rect 36180 15734 36210 16906
rect 36060 15720 36210 15734
rect 36270 15720 36360 16920
rect 36420 16906 36600 16920
rect 36420 15734 36450 16906
rect 36570 16320 36600 16906
rect 36660 16906 36810 16920
rect 36660 16334 36690 16906
rect 36660 16320 36810 16334
rect 37740 16906 37890 16920
rect 37860 16334 37890 16906
rect 37740 16320 37890 16334
rect 37950 16906 38130 16920
rect 37950 16334 37980 16906
rect 38100 16334 38130 16906
rect 37950 16320 38130 16334
rect 38190 16906 38340 16920
rect 38190 16334 38220 16906
rect 38190 16320 38340 16334
rect 38700 16906 38850 16920
rect 36420 15720 36570 15734
rect 38820 15734 38850 16906
rect 38700 15720 38850 15734
rect 38910 16860 39120 16920
rect 38910 15990 38954 16860
rect 39076 15990 39120 16860
rect 38910 15720 39120 15990
rect 39180 15720 39270 16920
rect 39330 16906 39630 16920
rect 39330 15734 39420 16906
rect 39540 15734 39630 16906
rect 39330 15720 39630 15734
rect 39690 15720 39780 16920
rect 39840 16860 40050 16920
rect 39840 15990 39884 16860
rect 40006 15990 40050 16860
rect 39840 15720 40050 15990
rect 40110 16906 40260 16920
rect 40110 15734 40140 16906
rect 40110 15720 40260 15734
rect 41580 16906 41730 16920
rect 41700 15734 41730 16906
rect 41580 15720 41730 15734
rect 41790 16860 42000 16920
rect 41790 15990 41834 16860
rect 41956 15990 42000 16860
rect 41790 15720 42000 15990
rect 42060 15720 42150 16920
rect 42210 16906 42510 16920
rect 42210 15734 42300 16906
rect 42420 15734 42510 16906
rect 42210 15720 42510 15734
rect 42570 15720 42660 16920
rect 42720 16860 42930 16920
rect 42720 15990 42764 16860
rect 42886 15990 42930 16860
rect 42720 15720 42930 15990
rect 42990 16906 43140 16920
rect 42990 15734 43020 16906
rect 42990 15720 43140 15734
rect 44460 16906 44610 16920
rect 44580 15734 44610 16906
rect 44460 15720 44610 15734
rect 44670 15720 44760 16920
rect 44820 16906 45000 16920
rect 44820 15734 44850 16906
rect 44970 16320 45000 16906
rect 45060 16906 45210 16920
rect 45060 16334 45090 16906
rect 45060 16320 45210 16334
rect 46140 16906 46290 16920
rect 46260 16334 46290 16906
rect 46140 16320 46290 16334
rect 46350 16906 46530 16920
rect 46350 16334 46380 16906
rect 46500 16334 46530 16906
rect 46350 16320 46530 16334
rect 46590 16906 46740 16920
rect 46590 16334 46620 16906
rect 46590 16320 46740 16334
rect 47580 16906 47730 16920
rect 47700 16334 47730 16906
rect 47580 16320 47730 16334
rect 47790 16906 47970 16920
rect 47790 16334 47820 16906
rect 47940 16334 47970 16906
rect 47790 16320 47970 16334
rect 48030 16906 48180 16920
rect 48030 16334 48060 16906
rect 48030 16320 48180 16334
rect 49020 16906 49170 16920
rect 44820 15720 44970 15734
rect 49140 15734 49170 16906
rect 49020 15720 49170 15734
rect 49230 15720 49320 16920
rect 49380 16906 49560 16920
rect 49380 15734 49410 16906
rect 49530 16320 49560 16906
rect 49620 16906 49770 16920
rect 49620 16334 49650 16906
rect 49620 16320 49770 16334
rect 49380 15720 49530 15734
rect 8940 12466 9090 12480
rect 6780 11866 6930 11880
rect 6900 11294 6930 11866
rect 6780 11280 6930 11294
rect 6990 11866 7170 11880
rect 6990 11294 7020 11866
rect 7140 11294 7170 11866
rect 6990 11280 7170 11294
rect 7230 11866 7380 11880
rect 7230 11294 7260 11866
rect 7230 11280 7380 11294
rect 9060 11294 9090 12466
rect 8940 11280 9090 11294
rect 9150 11280 9240 12480
rect 9300 12466 9660 12480
rect 9300 11294 9344 12466
rect 9616 11294 9660 12466
rect 9300 11280 9660 11294
rect 9720 11280 9810 12480
rect 9870 12466 10020 12480
rect 9870 11294 9900 12466
rect 12390 12466 12540 12480
rect 9870 11280 10020 11294
rect 10860 11866 11010 11880
rect 10980 11294 11010 11866
rect 10860 11280 11010 11294
rect 11070 11866 11250 11880
rect 11070 11294 11100 11866
rect 11220 11294 11250 11866
rect 11070 11280 11250 11294
rect 11310 11866 11460 11880
rect 11310 11294 11340 11866
rect 11310 11280 11460 11294
rect 12150 11866 12300 11880
rect 12270 11294 12300 11866
rect 12150 11280 12300 11294
rect 12360 11294 12390 11880
rect 12510 11294 12540 12466
rect 12360 11280 12540 11294
rect 12600 11280 12690 12480
rect 12750 12466 12900 12480
rect 12750 11294 12780 12466
rect 16950 12466 17100 12480
rect 12750 11280 12900 11294
rect 15900 11866 16050 11880
rect 16020 11294 16050 11866
rect 15900 11280 16050 11294
rect 16110 11866 16290 11880
rect 16110 11294 16140 11866
rect 16260 11294 16290 11866
rect 16110 11280 16290 11294
rect 16350 11866 16500 11880
rect 16350 11294 16380 11866
rect 16350 11280 16500 11294
rect 16710 11866 16860 11880
rect 16830 11294 16860 11866
rect 16710 11280 16860 11294
rect 16920 11294 16950 11880
rect 17070 11294 17100 12466
rect 16920 11280 17100 11294
rect 17160 11280 17250 12480
rect 17310 12466 17460 12480
rect 17310 11294 17340 12466
rect 17310 11280 17460 11294
rect 17580 12466 17730 12480
rect 17700 11294 17730 12466
rect 17580 11280 17730 11294
rect 17790 12210 18000 12480
rect 17790 11340 17834 12210
rect 17956 11340 18000 12210
rect 17790 11280 18000 11340
rect 18060 11280 18150 12480
rect 18210 12466 18510 12480
rect 18210 11294 18300 12466
rect 18420 11294 18510 12466
rect 18210 11280 18510 11294
rect 18570 11280 18660 12480
rect 18720 12210 18930 12480
rect 18720 11340 18764 12210
rect 18886 11340 18930 12210
rect 18720 11280 18930 11340
rect 18990 12466 19140 12480
rect 18990 11294 19020 12466
rect 18990 11280 19140 11294
rect 19260 12466 19410 12480
rect 19380 11294 19410 12466
rect 19260 11280 19410 11294
rect 19470 12210 19680 12480
rect 19470 11340 19514 12210
rect 19636 11340 19680 12210
rect 19470 11280 19680 11340
rect 19740 11280 19830 12480
rect 19890 12466 20190 12480
rect 19890 11294 19980 12466
rect 20100 11294 20190 12466
rect 19890 11280 20190 11294
rect 20250 11280 20340 12480
rect 20400 12210 20610 12480
rect 20400 11340 20444 12210
rect 20566 11340 20610 12210
rect 20400 11280 20610 11340
rect 20670 12466 20820 12480
rect 20670 11294 20700 12466
rect 20670 11280 20820 11294
rect 21900 12466 22050 12480
rect 22020 11294 22050 12466
rect 21900 11280 22050 11294
rect 22110 12210 22320 12480
rect 22110 11340 22154 12210
rect 22276 11340 22320 12210
rect 22110 11280 22320 11340
rect 22380 11280 22470 12480
rect 22530 12466 22830 12480
rect 22530 11294 22620 12466
rect 22740 11294 22830 12466
rect 22530 11280 22830 11294
rect 22890 11280 22980 12480
rect 23040 12210 23250 12480
rect 23040 11340 23084 12210
rect 23206 11340 23250 12210
rect 23040 11280 23250 11340
rect 23310 12466 23460 12480
rect 23310 11294 23340 12466
rect 23310 11280 23460 11294
rect 25020 12466 25170 12480
rect 25140 11294 25170 12466
rect 25020 11280 25170 11294
rect 25230 11280 25320 12480
rect 25380 12466 25530 12480
rect 25380 11294 25410 12466
rect 29100 12466 29250 12480
rect 25530 11294 25560 11880
rect 25380 11280 25560 11294
rect 25620 11866 25770 11880
rect 25620 11294 25650 11866
rect 25620 11280 25770 11294
rect 26700 11866 26850 11880
rect 26820 11294 26850 11866
rect 26700 11280 26850 11294
rect 26910 11866 27090 11880
rect 26910 11294 26940 11866
rect 27060 11294 27090 11866
rect 26910 11280 27090 11294
rect 27150 11866 27300 11880
rect 27150 11294 27180 11866
rect 27150 11280 27300 11294
rect 29220 11294 29250 12466
rect 29100 11280 29250 11294
rect 29310 11280 29400 12480
rect 29460 12466 29610 12480
rect 29460 11294 29490 12466
rect 30630 12466 30780 12480
rect 29610 11294 29640 11880
rect 29460 11280 29640 11294
rect 29700 11866 29850 11880
rect 29700 11294 29730 11866
rect 29700 11280 29850 11294
rect 30390 11866 30540 11880
rect 30510 11294 30540 11866
rect 30390 11280 30540 11294
rect 30600 11294 30630 11880
rect 30750 11294 30780 12466
rect 30600 11280 30780 11294
rect 30840 11280 30930 12480
rect 30990 12466 31140 12480
rect 30990 11294 31020 12466
rect 32940 12466 33090 12480
rect 30990 11280 31140 11294
rect 31980 11866 32130 11880
rect 32100 11294 32130 11866
rect 31980 11280 32130 11294
rect 32190 11866 32370 11880
rect 32190 11294 32220 11866
rect 32340 11294 32370 11866
rect 32190 11280 32370 11294
rect 32430 11866 32580 11880
rect 32430 11294 32460 11866
rect 32430 11280 32580 11294
rect 33060 11294 33090 12466
rect 32940 11280 33090 11294
rect 33150 12210 33360 12480
rect 33150 11340 33194 12210
rect 33316 11340 33360 12210
rect 33150 11280 33360 11340
rect 33420 11280 33510 12480
rect 33570 12466 33870 12480
rect 33570 11294 33660 12466
rect 33780 11294 33870 12466
rect 33570 11280 33870 11294
rect 33930 11280 34020 12480
rect 34080 12210 34290 12480
rect 34080 11340 34124 12210
rect 34246 11340 34290 12210
rect 34080 11280 34290 11340
rect 34350 12466 34500 12480
rect 34350 11294 34380 12466
rect 34350 11280 34500 11294
rect 34620 12466 34770 12480
rect 34740 11294 34770 12466
rect 34620 11280 34770 11294
rect 34830 11280 34920 12480
rect 34980 12466 35130 12480
rect 34980 11294 35010 12466
rect 40470 12466 40620 12480
rect 35130 11294 35160 11880
rect 34980 11280 35160 11294
rect 35220 11866 35370 11880
rect 35220 11294 35250 11866
rect 35220 11280 35370 11294
rect 36060 11866 36210 11880
rect 36180 11294 36210 11866
rect 36060 11280 36210 11294
rect 36270 11866 36450 11880
rect 36270 11294 36300 11866
rect 36420 11294 36450 11866
rect 36270 11280 36450 11294
rect 36510 11866 36660 11880
rect 36510 11294 36540 11866
rect 36510 11280 36660 11294
rect 37500 11866 37650 11880
rect 37620 11294 37650 11866
rect 37500 11280 37650 11294
rect 37710 11866 37890 11880
rect 37710 11294 37740 11866
rect 37860 11294 37890 11866
rect 37710 11280 37890 11294
rect 37950 11866 38100 11880
rect 37950 11294 37980 11866
rect 37950 11280 38100 11294
rect 38940 11866 39090 11880
rect 39060 11294 39090 11866
rect 38940 11280 39090 11294
rect 39150 11866 39330 11880
rect 39150 11294 39180 11866
rect 39300 11294 39330 11866
rect 39150 11280 39330 11294
rect 39390 11866 39540 11880
rect 39390 11294 39420 11866
rect 39390 11280 39540 11294
rect 40230 11866 40380 11880
rect 40350 11294 40380 11866
rect 40230 11280 40380 11294
rect 40440 11294 40470 11880
rect 40590 11294 40620 12466
rect 40440 11280 40620 11294
rect 40680 11280 40770 12480
rect 40830 12466 40980 12480
rect 40830 11294 40860 12466
rect 44460 12466 44610 12480
rect 40830 11280 40980 11294
rect 41580 11866 41730 11880
rect 41700 11294 41730 11866
rect 41580 11280 41730 11294
rect 41790 11866 41970 11880
rect 41790 11294 41820 11866
rect 41940 11294 41970 11866
rect 41790 11280 41970 11294
rect 42030 11866 42210 11880
rect 42030 11294 42060 11866
rect 42180 11294 42210 11866
rect 42030 11280 42210 11294
rect 42270 11866 42420 11880
rect 42270 11294 42300 11866
rect 42270 11280 42420 11294
rect 43260 11866 43410 11880
rect 43380 11294 43410 11866
rect 43260 11280 43410 11294
rect 43470 11866 43650 11880
rect 43470 11294 43500 11866
rect 43620 11294 43650 11866
rect 43470 11280 43650 11294
rect 43710 11866 43860 11880
rect 43710 11294 43740 11866
rect 43710 11280 43860 11294
rect 44580 11294 44610 12466
rect 44460 11280 44610 11294
rect 44670 11280 44760 12480
rect 44820 12466 44970 12480
rect 44820 11294 44850 12466
rect 47580 12466 47730 12480
rect 44970 11294 45000 11880
rect 44820 11280 45000 11294
rect 45060 11866 45210 11880
rect 45060 11294 45090 11866
rect 45060 11280 45210 11294
rect 46140 11866 46290 11880
rect 46260 11294 46290 11866
rect 46140 11280 46290 11294
rect 46350 11866 46530 11880
rect 46350 11294 46380 11866
rect 46500 11294 46530 11866
rect 46350 11280 46530 11294
rect 46590 11866 46740 11880
rect 46590 11294 46620 11866
rect 46590 11280 46740 11294
rect 47700 11294 47730 12466
rect 47580 11280 47730 11294
rect 47790 11280 47880 12480
rect 47940 12466 48090 12480
rect 47940 11294 47970 12466
rect 48090 11294 48120 11880
rect 47940 11280 48120 11294
rect 48180 11866 48330 11880
rect 48180 11294 48210 11866
rect 48180 11280 48330 11294
rect 49260 11866 49410 11880
rect 49380 11294 49410 11866
rect 49260 11280 49410 11294
rect 49470 11866 49650 11880
rect 49470 11294 49500 11866
rect 49620 11294 49650 11866
rect 49470 11280 49650 11294
rect 49710 11866 49860 11880
rect 49710 11294 49740 11866
rect 49710 11280 49860 11294
rect 5670 10906 5820 10920
rect 5790 10334 5820 10906
rect 5670 10320 5820 10334
rect 5880 10906 6060 10920
rect 5880 10320 5910 10906
rect 6030 9734 6060 10906
rect 5910 9720 6060 9734
rect 6120 9720 6210 10920
rect 6270 10906 6420 10920
rect 6270 9734 6300 10906
rect 6780 10906 6930 10920
rect 6900 10334 6930 10906
rect 6780 10320 6930 10334
rect 6990 10906 7170 10920
rect 6990 10334 7020 10906
rect 7140 10334 7170 10906
rect 6990 10320 7170 10334
rect 7230 10906 7380 10920
rect 7230 10334 7260 10906
rect 7230 10320 7380 10334
rect 7740 10906 7890 10920
rect 6270 9720 6420 9734
rect 7860 9734 7890 10906
rect 7740 9720 7890 9734
rect 7950 10860 8160 10920
rect 7950 9990 7994 10860
rect 8116 9990 8160 10860
rect 7950 9720 8160 9990
rect 8220 9720 8310 10920
rect 8370 10906 8670 10920
rect 8370 9734 8460 10906
rect 8580 9734 8670 10906
rect 8370 9720 8670 9734
rect 8730 9720 8820 10920
rect 8880 10860 9090 10920
rect 8880 9990 8924 10860
rect 9046 9990 9090 10860
rect 8880 9720 9090 9990
rect 9150 10906 9300 10920
rect 9150 9734 9180 10906
rect 9660 10906 9810 10920
rect 9780 10334 9810 10906
rect 9660 10320 9810 10334
rect 9870 10906 10050 10920
rect 9870 10334 9900 10906
rect 10020 10334 10050 10906
rect 9870 10320 10050 10334
rect 10110 10906 10290 10920
rect 10110 10334 10140 10906
rect 10260 10334 10290 10906
rect 10110 10320 10290 10334
rect 10350 10906 10500 10920
rect 10350 10334 10380 10906
rect 10350 10320 10500 10334
rect 11340 10906 11490 10920
rect 11460 10334 11490 10906
rect 11340 10320 11490 10334
rect 11550 10906 11730 10920
rect 11550 10334 11580 10906
rect 11700 10334 11730 10906
rect 11550 10320 11730 10334
rect 11790 10906 11940 10920
rect 11790 10334 11820 10906
rect 11790 10320 11940 10334
rect 13740 10906 13890 10920
rect 9150 9720 9300 9734
rect 13860 9734 13890 10906
rect 13740 9720 13890 9734
rect 13950 10860 14160 10920
rect 13950 9990 13994 10860
rect 14116 9990 14160 10860
rect 13950 9720 14160 9990
rect 14220 9720 14310 10920
rect 14370 10906 14670 10920
rect 14370 9734 14460 10906
rect 14580 9734 14670 10906
rect 14370 9720 14670 9734
rect 14730 9720 14820 10920
rect 14880 10860 15090 10920
rect 14880 9990 14924 10860
rect 15046 9990 15090 10860
rect 14880 9720 15090 9990
rect 15150 10906 15300 10920
rect 15150 9734 15180 10906
rect 16380 10906 16530 10920
rect 16500 10334 16530 10906
rect 16380 10320 16530 10334
rect 16590 10906 16770 10920
rect 16590 10334 16620 10906
rect 16740 10334 16770 10906
rect 16590 10320 16770 10334
rect 16830 10906 16980 10920
rect 16830 10334 16860 10906
rect 16830 10320 16980 10334
rect 17340 10906 17490 10920
rect 15150 9720 15300 9734
rect 17460 9734 17490 10906
rect 17340 9720 17490 9734
rect 17550 10860 17760 10920
rect 17550 9990 17594 10860
rect 17716 9990 17760 10860
rect 17550 9720 17760 9990
rect 17820 9720 17910 10920
rect 17970 10906 18270 10920
rect 17970 9734 18060 10906
rect 18180 9734 18270 10906
rect 17970 9720 18270 9734
rect 18330 9720 18420 10920
rect 18480 10860 18690 10920
rect 18480 9990 18524 10860
rect 18646 9990 18690 10860
rect 18480 9720 18690 9990
rect 18750 10906 18900 10920
rect 18750 9734 18780 10906
rect 18750 9720 18900 9734
rect 19260 10906 19410 10920
rect 19380 9734 19410 10906
rect 19260 9720 19410 9734
rect 19470 10860 19680 10920
rect 19470 9990 19514 10860
rect 19636 9990 19680 10860
rect 19470 9720 19680 9990
rect 19740 9720 19830 10920
rect 19890 10906 20190 10920
rect 19890 9734 19980 10906
rect 20100 9734 20190 10906
rect 19890 9720 20190 9734
rect 20250 9720 20340 10920
rect 20400 10860 20610 10920
rect 20400 9990 20444 10860
rect 20566 9990 20610 10860
rect 20400 9720 20610 9990
rect 20670 10906 20820 10920
rect 20670 9734 20700 10906
rect 21180 10906 21330 10920
rect 21300 10334 21330 10906
rect 21180 10320 21330 10334
rect 21390 10906 21570 10920
rect 21390 10334 21420 10906
rect 21540 10334 21570 10906
rect 21390 10320 21570 10334
rect 21630 10906 21780 10920
rect 21630 10334 21660 10906
rect 21630 10320 21780 10334
rect 21900 10906 22050 10920
rect 20670 9720 20820 9734
rect 22020 9734 22050 10906
rect 21900 9720 22050 9734
rect 22110 10860 22320 10920
rect 22110 9990 22154 10860
rect 22276 9990 22320 10860
rect 22110 9720 22320 9990
rect 22380 9720 22470 10920
rect 22530 10906 22830 10920
rect 22530 9734 22620 10906
rect 22740 9734 22830 10906
rect 22530 9720 22830 9734
rect 22890 9720 22980 10920
rect 23040 10860 23250 10920
rect 23040 9990 23084 10860
rect 23206 9990 23250 10860
rect 23040 9720 23250 9990
rect 23310 10906 23460 10920
rect 23310 9734 23340 10906
rect 23820 10906 23970 10920
rect 23940 10334 23970 10906
rect 23820 10320 23970 10334
rect 24030 10906 24210 10920
rect 24030 10334 24060 10906
rect 24180 10334 24210 10906
rect 24030 10320 24210 10334
rect 24270 10906 24420 10920
rect 24270 10334 24300 10906
rect 24270 10320 24420 10334
rect 25500 10906 25650 10920
rect 23310 9720 23460 9734
rect 25620 9734 25650 10906
rect 25500 9720 25650 9734
rect 25710 10860 25920 10920
rect 25710 9990 25754 10860
rect 25876 9990 25920 10860
rect 25710 9720 25920 9990
rect 25980 9720 26070 10920
rect 26130 10906 26430 10920
rect 26130 9734 26220 10906
rect 26340 9734 26430 10906
rect 26130 9720 26430 9734
rect 26490 9720 26580 10920
rect 26640 10860 26850 10920
rect 26640 9990 26684 10860
rect 26806 9990 26850 10860
rect 26640 9720 26850 9990
rect 26910 10906 27060 10920
rect 26910 9734 26940 10906
rect 27900 10906 28050 10920
rect 28020 10334 28050 10906
rect 27900 10320 28050 10334
rect 28110 10906 28290 10920
rect 28110 10334 28140 10906
rect 28260 10334 28290 10906
rect 28110 10320 28290 10334
rect 28350 10906 28500 10920
rect 28350 10334 28380 10906
rect 28350 10320 28500 10334
rect 29340 10890 29490 10920
rect 29460 10320 29490 10890
rect 29550 10890 29700 10920
rect 29550 10320 29580 10890
rect 30540 10890 30690 10920
rect 30660 10320 30690 10890
rect 30750 10890 30900 10920
rect 30750 10320 30780 10890
rect 31740 10906 31890 10920
rect 26910 9720 27060 9734
rect 31860 9734 31890 10906
rect 31740 9720 31890 9734
rect 31950 9720 32040 10920
rect 32100 10906 32280 10920
rect 32100 9734 32130 10906
rect 32250 10320 32280 10906
rect 32340 10906 32490 10920
rect 32340 10334 32370 10906
rect 32340 10320 32490 10334
rect 33180 10906 33330 10920
rect 32100 9720 32250 9734
rect 33300 9734 33330 10906
rect 33180 9720 33330 9734
rect 33390 10860 33600 10920
rect 33390 9990 33434 10860
rect 33556 9990 33600 10860
rect 33390 9720 33600 9990
rect 33660 9720 33750 10920
rect 33810 10906 34110 10920
rect 33810 9734 33900 10906
rect 34020 9734 34110 10906
rect 33810 9720 34110 9734
rect 34170 9720 34260 10920
rect 34320 10860 34530 10920
rect 34320 9990 34364 10860
rect 34486 9990 34530 10860
rect 34320 9720 34530 9990
rect 34590 10906 34740 10920
rect 34590 9734 34620 10906
rect 35580 10906 35730 10920
rect 35700 10334 35730 10906
rect 35580 10320 35730 10334
rect 35790 10906 35970 10920
rect 35790 10334 35820 10906
rect 35940 10334 35970 10906
rect 35790 10320 35970 10334
rect 36030 10906 36210 10920
rect 36030 10334 36060 10906
rect 36180 10334 36210 10906
rect 36030 10320 36210 10334
rect 36270 10906 36420 10920
rect 36270 10334 36300 10906
rect 36270 10320 36420 10334
rect 36780 10906 36930 10920
rect 36900 10334 36930 10906
rect 36780 10320 36930 10334
rect 36990 10906 37170 10920
rect 36990 10334 37020 10906
rect 37140 10334 37170 10906
rect 36990 10320 37170 10334
rect 37230 10906 37380 10920
rect 37230 10334 37260 10906
rect 37230 10320 37380 10334
rect 37740 10906 37890 10920
rect 37860 10334 37890 10906
rect 37740 10320 37890 10334
rect 37950 10906 38130 10920
rect 37950 10334 37980 10906
rect 38100 10334 38130 10906
rect 37950 10320 38130 10334
rect 38190 10906 38370 10920
rect 38190 10334 38220 10906
rect 38340 10334 38370 10906
rect 38190 10320 38370 10334
rect 38430 10906 38580 10920
rect 38430 10334 38460 10906
rect 38430 10320 38580 10334
rect 38940 10906 39090 10920
rect 34590 9720 34740 9734
rect 39060 9734 39090 10906
rect 38940 9720 39090 9734
rect 39150 9720 39240 10920
rect 39300 10906 39480 10920
rect 39300 9734 39330 10906
rect 39450 10320 39480 10906
rect 39540 10906 39690 10920
rect 39540 10334 39570 10906
rect 39540 10320 39690 10334
rect 40380 10906 40530 10920
rect 40500 10334 40530 10906
rect 40380 10320 40530 10334
rect 40590 10906 40770 10920
rect 40590 10334 40620 10906
rect 40740 10334 40770 10906
rect 40590 10320 40770 10334
rect 40830 10906 40980 10920
rect 40830 10334 40860 10906
rect 40830 10320 40980 10334
rect 41580 10906 41730 10920
rect 41700 10334 41730 10906
rect 41580 10320 41730 10334
rect 41790 10906 41970 10920
rect 41790 10334 41820 10906
rect 41940 10334 41970 10906
rect 41790 10320 41970 10334
rect 42030 10906 42180 10920
rect 42030 10334 42060 10906
rect 42030 10320 42180 10334
rect 42540 10906 42690 10920
rect 39300 9720 39450 9734
rect 42660 9734 42690 10906
rect 42540 9720 42690 9734
rect 42750 10860 42960 10920
rect 42750 9990 42794 10860
rect 42916 9990 42960 10860
rect 42750 9720 42960 9990
rect 43020 9720 43110 10920
rect 43170 10906 43470 10920
rect 43170 9734 43260 10906
rect 43380 9734 43470 10906
rect 43170 9720 43470 9734
rect 43530 9720 43620 10920
rect 43680 10860 43890 10920
rect 43680 9990 43724 10860
rect 43846 9990 43890 10860
rect 43680 9720 43890 9990
rect 43950 10906 44100 10920
rect 43950 9734 43980 10906
rect 43950 9720 44100 9734
rect 45180 10906 45330 10920
rect 45300 9734 45330 10906
rect 45180 9720 45330 9734
rect 45390 10860 45600 10920
rect 45390 9990 45434 10860
rect 45556 9990 45600 10860
rect 45390 9720 45600 9990
rect 45660 9720 45750 10920
rect 45810 10906 46110 10920
rect 45810 9734 45900 10906
rect 46020 9734 46110 10906
rect 45810 9720 46110 9734
rect 46170 9720 46260 10920
rect 46320 10860 46530 10920
rect 46320 9990 46364 10860
rect 46486 9990 46530 10860
rect 46320 9720 46530 9990
rect 46590 10906 46740 10920
rect 46590 9734 46620 10906
rect 47580 10906 47730 10920
rect 47700 10334 47730 10906
rect 47580 10320 47730 10334
rect 47790 10906 47970 10920
rect 47790 10334 47820 10906
rect 47940 10334 47970 10906
rect 47790 10320 47970 10334
rect 48030 10906 48180 10920
rect 48030 10334 48060 10906
rect 48030 10320 48180 10334
rect 49020 10906 49170 10920
rect 49140 10334 49170 10906
rect 49020 10320 49170 10334
rect 49230 10906 49410 10920
rect 49230 10334 49260 10906
rect 49380 10334 49410 10906
rect 49230 10320 49410 10334
rect 49470 10906 49620 10920
rect 49470 10334 49500 10906
rect 49470 10320 49620 10334
rect 46590 9720 46740 9734
rect 5580 6466 5730 6480
rect 5700 5294 5730 6466
rect 5580 5280 5730 5294
rect 5790 6210 6000 6480
rect 5790 5340 5834 6210
rect 5956 5340 6000 6210
rect 5790 5280 6000 5340
rect 6060 5280 6150 6480
rect 6210 6466 6510 6480
rect 6210 5294 6300 6466
rect 6420 5294 6510 6466
rect 6210 5280 6510 5294
rect 6570 5280 6660 6480
rect 6720 6210 6930 6480
rect 6720 5340 6764 6210
rect 6886 5340 6930 6210
rect 6720 5280 6930 5340
rect 6990 6466 7140 6480
rect 6990 5294 7020 6466
rect 9030 6466 9180 6480
rect 6990 5280 7140 5294
rect 8100 5310 8130 5880
rect 7980 5280 8130 5310
rect 8190 5310 8220 5880
rect 8190 5280 8340 5310
rect 8790 5866 8940 5880
rect 8910 5294 8940 5866
rect 8790 5280 8940 5294
rect 9000 5294 9030 5880
rect 9150 5294 9180 6466
rect 9000 5280 9180 5294
rect 9240 5280 9330 6480
rect 9390 6466 9540 6480
rect 9390 5294 9420 6466
rect 11190 6466 11340 6480
rect 9390 5280 9540 5294
rect 9900 5866 10050 5880
rect 10020 5294 10050 5866
rect 9900 5280 10050 5294
rect 10110 5866 10290 5880
rect 10110 5294 10140 5866
rect 10260 5294 10290 5866
rect 10110 5280 10290 5294
rect 10350 5866 10500 5880
rect 10350 5294 10380 5866
rect 10350 5280 10500 5294
rect 10950 5866 11100 5880
rect 11070 5294 11100 5866
rect 10950 5280 11100 5294
rect 11160 5294 11190 5880
rect 11310 5294 11340 6466
rect 11160 5280 11340 5294
rect 11400 5280 11490 6480
rect 11550 6466 11700 6480
rect 11550 5294 11580 6466
rect 13740 6346 13890 6480
rect 11550 5280 11700 5294
rect 12300 5866 12450 5880
rect 12420 5294 12450 5866
rect 12300 5280 12450 5294
rect 12510 5866 12690 5880
rect 12510 5294 12540 5866
rect 12660 5294 12690 5866
rect 12510 5280 12690 5294
rect 12750 5866 12900 5880
rect 12750 5294 12780 5866
rect 12750 5280 12900 5294
rect 13860 5324 13890 6346
rect 13740 5280 13890 5324
rect 13950 6300 14130 6480
rect 13950 5280 13980 6300
rect 14100 5280 14130 6300
rect 14190 6466 14370 6480
rect 14190 5294 14220 6466
rect 14340 5294 14370 6466
rect 14190 5280 14370 5294
rect 14430 6466 14580 6480
rect 14430 5294 14460 6466
rect 14430 5280 14580 5294
rect 15540 5310 15570 6480
rect 15420 5280 15570 5310
rect 15630 5280 15720 6480
rect 15780 5310 15810 6480
rect 15780 5280 15930 5310
rect 18180 5310 18210 6480
rect 18060 5280 18210 5310
rect 18270 5280 18360 6480
rect 18420 5310 18450 6480
rect 25740 6466 25890 6480
rect 18420 5280 18570 5310
rect 20700 5866 20850 5880
rect 20820 5294 20850 5866
rect 20700 5280 20850 5294
rect 20910 5866 21090 5880
rect 20910 5294 20940 5866
rect 21060 5294 21090 5866
rect 20910 5280 21090 5294
rect 21150 5866 21300 5880
rect 21150 5294 21180 5866
rect 21150 5280 21300 5294
rect 23340 5866 23490 5880
rect 23460 5294 23490 5866
rect 23340 5280 23490 5294
rect 23550 5866 23730 5880
rect 23550 5294 23580 5866
rect 23700 5294 23730 5866
rect 23550 5280 23730 5294
rect 23790 5866 23940 5880
rect 23790 5294 23820 5866
rect 23790 5280 23940 5294
rect 25860 5294 25890 6466
rect 25740 5280 25890 5294
rect 25950 6210 26160 6480
rect 25950 5340 25994 6210
rect 26116 5340 26160 6210
rect 25950 5280 26160 5340
rect 26220 5280 26310 6480
rect 26370 6466 26670 6480
rect 26370 5294 26460 6466
rect 26580 5294 26670 6466
rect 26370 5280 26670 5294
rect 26730 5280 26820 6480
rect 26880 6210 27090 6480
rect 26880 5340 26924 6210
rect 27046 5340 27090 6210
rect 26880 5280 27090 5340
rect 27150 6466 27300 6480
rect 27150 5294 27180 6466
rect 30060 6466 30210 6480
rect 27150 5280 27300 5294
rect 27900 5866 28050 5880
rect 28020 5294 28050 5866
rect 27900 5280 28050 5294
rect 28110 5866 28290 5880
rect 28110 5294 28140 5866
rect 28260 5294 28290 5866
rect 28110 5280 28290 5294
rect 28350 5866 28500 5880
rect 28350 5294 28380 5866
rect 28350 5280 28500 5294
rect 29100 5866 29250 5880
rect 29220 5294 29250 5866
rect 29100 5280 29250 5294
rect 29310 5866 29490 5880
rect 29310 5294 29340 5866
rect 29460 5294 29490 5866
rect 29310 5280 29490 5294
rect 29550 5866 29700 5880
rect 29550 5294 29580 5866
rect 29550 5280 29700 5294
rect 30180 5294 30210 6466
rect 30060 5280 30210 5294
rect 30270 6210 30480 6480
rect 30270 5340 30314 6210
rect 30436 5340 30480 6210
rect 30270 5280 30480 5340
rect 30540 5280 30630 6480
rect 30690 6466 30990 6480
rect 30690 5294 30780 6466
rect 30900 5294 30990 6466
rect 30690 5280 30990 5294
rect 31050 5280 31140 6480
rect 31200 6210 31410 6480
rect 31200 5340 31244 6210
rect 31366 5340 31410 6210
rect 31200 5280 31410 5340
rect 31470 6466 31620 6480
rect 31470 5294 31500 6466
rect 31470 5280 31620 5294
rect 31980 6466 32130 6480
rect 32100 5294 32130 6466
rect 31980 5280 32130 5294
rect 32190 5280 32280 6480
rect 32340 6466 32490 6480
rect 32340 5294 32370 6466
rect 37830 6466 37980 6480
rect 32490 5294 32520 5880
rect 32340 5280 32520 5294
rect 32580 5866 32730 5880
rect 32580 5294 32610 5866
rect 32580 5280 32730 5294
rect 33180 5866 33330 5880
rect 33300 5294 33330 5866
rect 33180 5280 33330 5294
rect 33390 5866 33570 5880
rect 33390 5294 33420 5866
rect 33540 5294 33570 5866
rect 33390 5280 33570 5294
rect 33630 5866 33780 5880
rect 33630 5294 33660 5866
rect 33630 5280 33780 5294
rect 34620 5866 34770 5880
rect 34740 5294 34770 5866
rect 34620 5280 34770 5294
rect 34830 5866 35010 5880
rect 34830 5294 34860 5866
rect 34980 5294 35010 5866
rect 34830 5280 35010 5294
rect 35070 5866 35220 5880
rect 35070 5294 35100 5866
rect 35070 5280 35220 5294
rect 36060 5866 36210 5880
rect 36180 5294 36210 5866
rect 36060 5280 36210 5294
rect 36270 5866 36450 5880
rect 36270 5294 36300 5866
rect 36420 5294 36450 5866
rect 36270 5280 36450 5294
rect 36510 5866 36660 5880
rect 36510 5294 36540 5866
rect 36510 5280 36660 5294
rect 37590 5866 37740 5880
rect 37710 5294 37740 5866
rect 37590 5280 37740 5294
rect 37800 5294 37830 5880
rect 37950 5294 37980 6466
rect 37800 5280 37980 5294
rect 38040 5280 38130 6480
rect 38190 6466 38340 6480
rect 38190 5294 38220 6466
rect 38190 5280 38340 5294
rect 38940 5866 39090 5880
rect 39060 5294 39090 5866
rect 38940 5280 39090 5294
rect 39150 5866 39330 5880
rect 39150 5294 39180 5866
rect 39300 5294 39330 5866
rect 39150 5280 39330 5294
rect 39390 5866 39540 5880
rect 39390 5294 39420 5866
rect 39390 5280 39540 5294
rect 40380 5866 40530 5880
rect 40500 5294 40530 5866
rect 40380 5280 40530 5294
rect 40590 5866 40770 5880
rect 40590 5294 40620 5866
rect 40740 5294 40770 5866
rect 40590 5280 40770 5294
rect 40830 5866 40980 5880
rect 40830 5294 40860 5866
rect 40830 5280 40980 5294
rect 43380 5310 43410 6480
rect 43260 5280 43410 5310
rect 43470 5280 43560 6480
rect 43620 5310 43650 6480
rect 43620 5280 43770 5310
rect 44460 6346 44610 6480
rect 44580 5324 44610 6346
rect 44460 5280 44610 5324
rect 44670 6300 44850 6480
rect 44670 5280 44700 6300
rect 44820 5280 44850 6300
rect 44910 6466 45090 6480
rect 44910 5294 44940 6466
rect 45060 5294 45090 6466
rect 44910 5280 45090 5294
rect 45150 5460 45180 6480
rect 45300 5460 45330 6480
rect 45150 5280 45330 5460
rect 45390 6466 45540 6480
rect 45390 5294 45420 6466
rect 47670 6466 47820 6480
rect 45390 5280 45540 5294
rect 46500 5310 46530 5880
rect 46380 5280 46530 5310
rect 46590 5310 46620 5880
rect 46590 5280 46740 5310
rect 47430 5866 47580 5880
rect 47550 5294 47580 5866
rect 47430 5280 47580 5294
rect 47640 5294 47670 5880
rect 47790 5294 47820 6466
rect 47640 5280 47820 5294
rect 47880 5280 47970 6480
rect 48030 6466 48180 6480
rect 48030 5294 48060 6466
rect 48030 5280 48180 5294
<< ndcontact >>
rect 5580 43320 5700 43920
rect 5820 43320 5940 43920
rect 6060 43470 6180 43890
rect 6300 43320 6420 43920
rect 6780 43320 6900 43920
rect 7170 43320 7290 43920
rect 7740 43320 7860 43920
rect 7980 43320 8100 43920
rect 8220 43470 8340 43890
rect 8460 43320 8580 43920
rect 8940 43320 9060 43920
rect 9180 43440 9330 43890
rect 9660 43440 9780 43860
rect 10110 43440 10260 43890
rect 10380 43320 10500 43920
rect 10860 43620 10980 43920
rect 11100 43620 11220 43920
rect 11340 43620 11460 43920
rect 12300 43620 12420 43920
rect 12540 43620 12660 43920
rect 12780 43620 12900 43920
rect 13740 43320 13860 43920
rect 13980 43470 14100 43890
rect 14220 43320 14340 43920
rect 14460 43320 14580 43920
rect 15420 43320 15540 43920
rect 15810 43320 15930 43920
rect 17100 43320 17220 43920
rect 17340 43470 17460 43890
rect 17580 43320 17700 43920
rect 17820 43320 17940 43920
rect 19260 43320 19380 43920
rect 19500 43440 19650 43890
rect 19980 43440 20100 43860
rect 20430 43440 20580 43890
rect 20700 43320 20820 43920
rect 21180 43650 21300 43920
rect 21420 43650 21540 43920
rect 22620 43320 22740 43920
rect 22860 43440 23010 43890
rect 23340 43440 23460 43860
rect 23790 43440 23940 43890
rect 24060 43320 24180 43920
rect 25020 43320 25140 43920
rect 25260 43320 25380 43920
rect 25500 43470 25620 43890
rect 25740 43320 25860 43920
rect 26700 43320 26820 43920
rect 27090 43320 27210 43920
rect 27900 43320 28020 43920
rect 28140 43470 28260 43890
rect 28380 43320 28500 43920
rect 28620 43320 28740 43920
rect 29100 43320 29220 43920
rect 29490 43320 29610 43920
rect 30300 43320 30420 43920
rect 30540 43470 30660 43890
rect 30780 43320 30900 43920
rect 31020 43320 31140 43920
rect 31740 43320 31860 43920
rect 31980 43470 32100 43890
rect 32220 43320 32340 43920
rect 32460 43320 32580 43920
rect 33270 43320 33390 43920
rect 33660 43320 33780 43920
rect 34620 43620 34740 43920
rect 34860 43620 34980 43920
rect 35100 43620 35220 43920
rect 35820 43320 35940 43920
rect 36060 43440 36210 43890
rect 36540 43440 36660 43860
rect 36990 43440 37140 43890
rect 37260 43320 37380 43920
rect 37740 43320 37860 43920
rect 37980 43320 38100 43920
rect 38220 43470 38340 43890
rect 38460 43320 38580 43920
rect 39420 43320 39540 43920
rect 39660 43440 39810 43890
rect 40140 43440 40260 43860
rect 40590 43440 40740 43890
rect 40860 43320 40980 43920
rect 41820 43650 41940 43920
rect 42060 43650 42180 43920
rect 43020 43320 43140 43920
rect 43260 43470 43380 43890
rect 43500 43320 43620 43920
rect 43740 43320 43860 43920
rect 44220 43320 44340 43920
rect 44460 43470 44580 43890
rect 44700 43320 44820 43920
rect 44940 43320 45060 43920
rect 45180 43650 45300 43920
rect 45420 43650 45540 43920
rect 45660 43320 45780 43920
rect 45900 43440 46050 43890
rect 46380 43440 46500 43860
rect 46830 43440 46980 43890
rect 47100 43320 47220 43920
rect 47340 43320 47460 43920
rect 47580 43440 47730 43890
rect 48060 43440 48180 43860
rect 48510 43440 48660 43890
rect 48780 43320 48900 43920
rect 5910 38280 6030 38880
rect 6300 38280 6420 38880
rect 6540 38280 6660 38580
rect 8310 38280 8430 38880
rect 8700 38280 8820 38880
rect 9660 38280 9780 38880
rect 10050 38280 10170 38880
rect 10620 38280 10740 38580
rect 10860 38280 10980 38880
rect 11250 38280 11370 38880
rect 11580 38280 11700 38880
rect 11820 38310 11970 38760
rect 12300 38340 12420 38760
rect 12750 38310 12900 38760
rect 13020 38280 13140 38880
rect 13500 38280 13620 38880
rect 13890 38280 14010 38880
rect 14550 38280 14670 38580
rect 14790 38280 14910 38880
rect 15180 38280 15300 38880
rect 15660 38280 15780 38550
rect 15900 38280 16020 38550
rect 16380 38280 16500 38880
rect 16620 38310 16740 38730
rect 16860 38280 16980 38880
rect 17100 38280 17220 38880
rect 17580 38280 17700 38880
rect 17820 38280 17940 38880
rect 18060 38310 18180 38730
rect 18300 38280 18420 38880
rect 18540 38280 18660 38550
rect 18780 38280 18900 38550
rect 19260 38280 19380 38880
rect 19500 38310 19620 38730
rect 19740 38280 19860 38880
rect 19980 38280 20100 38880
rect 21030 38280 21150 38880
rect 21420 38280 21540 38880
rect 21900 38280 22020 38880
rect 22140 38310 22290 38760
rect 22620 38340 22740 38760
rect 23070 38310 23220 38760
rect 23340 38280 23460 38880
rect 23820 38280 23940 38580
rect 24060 38280 24180 38580
rect 24300 38280 24420 38580
rect 24780 38280 24900 38880
rect 25020 38310 25140 38730
rect 25260 38280 25380 38880
rect 25500 38280 25620 38880
rect 26280 38280 26400 38880
rect 26730 38280 26850 38880
rect 27180 38280 27300 38880
rect 27900 38280 28020 38550
rect 28140 38280 28260 38550
rect 30630 38280 30750 38880
rect 31020 38280 31140 38880
rect 32070 38280 32190 38880
rect 32460 38280 32580 38880
rect 33420 38280 33540 38880
rect 33660 38310 33810 38760
rect 34140 38340 34260 38760
rect 34590 38310 34740 38760
rect 34860 38280 34980 38880
rect 36060 38280 36180 38880
rect 36300 38310 36420 38730
rect 36540 38280 36660 38880
rect 36780 38280 36900 38880
rect 37830 38280 37950 38880
rect 38220 38280 38340 38880
rect 38940 38280 39060 38880
rect 39180 38310 39300 38730
rect 39420 38280 39540 38880
rect 39660 38280 39780 38880
rect 40380 38280 40500 38880
rect 40770 38280 40890 38880
rect 41820 38280 41940 38550
rect 42060 38280 42180 38550
rect 43020 38280 43140 38880
rect 43260 38310 43380 38730
rect 43500 38280 43620 38880
rect 43740 38280 43860 38880
rect 44700 38280 44820 38550
rect 44940 38280 45060 38550
rect 45900 38280 46020 38880
rect 46140 38280 46260 38880
rect 46380 38310 46500 38730
rect 46620 38280 46740 38880
rect 47580 38280 47700 38880
rect 47820 38310 47940 38730
rect 48060 38280 48180 38880
rect 48300 38280 48420 38880
rect 49350 38280 49470 38880
rect 49740 38280 49860 38880
rect 5670 37320 5790 37920
rect 6060 37320 6180 37920
rect 7020 37740 7140 37890
rect 7260 37650 7380 37920
rect 8220 37320 8340 37920
rect 8460 37320 8580 37920
rect 8700 37470 8820 37890
rect 8940 37320 9060 37920
rect 10860 37320 10980 37920
rect 11250 37320 11370 37920
rect 12060 37320 12180 37920
rect 12300 37320 12420 37920
rect 12540 37470 12660 37890
rect 12780 37320 12900 37920
rect 14940 37320 15060 37920
rect 15180 37320 15300 37920
rect 15420 37470 15540 37890
rect 15660 37320 15780 37920
rect 16710 37620 16830 37920
rect 16950 37320 17070 37920
rect 17340 37320 17460 37920
rect 18060 37320 18180 37920
rect 18450 37320 18570 37920
rect 19500 37320 19620 37920
rect 19890 37320 20010 37920
rect 20940 37320 21060 37920
rect 21330 37320 21450 37920
rect 22380 37320 22500 37920
rect 22770 37320 22890 37920
rect 23820 37650 23940 37920
rect 24060 37650 24180 37920
rect 25110 37320 25230 37920
rect 25500 37320 25620 37920
rect 26460 37320 26580 37920
rect 26700 37470 26820 37890
rect 26940 37320 27060 37920
rect 27180 37320 27300 37920
rect 27900 37320 28020 37920
rect 28290 37320 28410 37920
rect 29100 37320 29220 37920
rect 29490 37320 29610 37920
rect 30060 37320 30180 37920
rect 30300 37470 30420 37890
rect 30540 37320 30660 37920
rect 30780 37320 30900 37920
rect 31260 37650 31380 37920
rect 31500 37650 31620 37920
rect 31980 37320 32100 37920
rect 32220 37320 32340 37920
rect 32460 37470 32580 37890
rect 32700 37320 32820 37920
rect 33270 37320 33390 37920
rect 33660 37320 33780 37920
rect 34620 37320 34740 37920
rect 35010 37320 35130 37920
rect 35580 37320 35700 37920
rect 35820 37440 35970 37890
rect 36300 37440 36420 37860
rect 36750 37440 36900 37890
rect 37020 37320 37140 37920
rect 38940 37650 39060 37920
rect 39180 37650 39300 37920
rect 39900 37320 40020 37920
rect 40350 37746 40470 37868
rect 40350 37402 40470 37522
rect 40800 37334 40920 37906
rect 41580 37650 41700 37920
rect 41820 37650 41940 37920
rect 42300 37334 42420 37906
rect 42540 37334 42660 37906
rect 42780 37470 42900 37890
rect 43020 37334 43140 37906
rect 43500 37650 43620 37920
rect 43740 37650 43860 37920
rect 44460 37334 44580 37906
rect 44700 37470 44820 37890
rect 44940 37334 45060 37906
rect 45180 37334 45300 37906
rect 46140 37334 46260 37906
rect 46530 37334 46650 37906
rect 47580 37334 47700 37906
rect 47820 37470 47940 37890
rect 48060 37334 48180 37906
rect 48300 37334 48420 37906
rect 49350 37334 49470 37906
rect 49740 37334 49860 37906
rect 6540 32294 6660 32866
rect 6780 32294 6900 32866
rect 7020 32310 7140 32730
rect 7260 32294 7380 32866
rect 7740 32294 7860 32866
rect 7980 32294 8100 32866
rect 8220 32310 8340 32730
rect 8460 32294 8580 32866
rect 8940 32294 9060 32866
rect 9194 32324 9316 32746
rect 9660 32340 9780 32760
rect 10124 32324 10246 32746
rect 10380 32294 10500 32866
rect 11100 32294 11220 32866
rect 11354 32324 11476 32746
rect 11820 32340 11940 32760
rect 12284 32324 12406 32746
rect 12540 32294 12660 32866
rect 13740 32280 13860 32550
rect 13980 32280 14100 32550
rect 15180 32294 15300 32866
rect 15570 32294 15690 32866
rect 16620 32294 16740 32866
rect 16860 32310 16980 32730
rect 17100 32294 17220 32866
rect 17340 32294 17460 32866
rect 19350 32294 19470 32866
rect 19740 32294 19860 32866
rect 20790 32294 20910 32566
rect 21030 32294 21150 32866
rect 21420 32294 21540 32866
rect 23340 32294 23460 32866
rect 23580 32310 23700 32730
rect 23820 32294 23940 32866
rect 24060 32294 24180 32866
rect 24780 32294 24900 32866
rect 25020 32310 25140 32730
rect 25260 32294 25380 32866
rect 25500 32294 25620 32866
rect 25980 32294 26100 32866
rect 26234 32324 26356 32746
rect 26700 32340 26820 32760
rect 27164 32324 27286 32746
rect 27420 32294 27540 32866
rect 30300 32280 30420 32550
rect 30540 32280 30660 32550
rect 31110 32294 31230 32866
rect 31500 32294 31620 32866
rect 31980 32294 32100 32866
rect 32220 32310 32340 32730
rect 32460 32294 32580 32866
rect 32700 32294 32820 32866
rect 33180 32294 33300 32866
rect 33570 32294 33690 32866
rect 34620 32294 34740 32866
rect 35010 32294 35130 32866
rect 36060 32294 36180 32866
rect 36450 32294 36570 32866
rect 37590 32294 37710 32866
rect 37980 32294 38100 32866
rect 38940 32294 39060 32866
rect 39330 32294 39450 32866
rect 40140 32294 40260 32866
rect 40380 32310 40500 32730
rect 40620 32294 40740 32866
rect 40860 32294 40980 32866
rect 41580 32294 41700 32866
rect 41970 32294 42090 32866
rect 43020 32294 43140 32866
rect 43260 32310 43380 32730
rect 43500 32294 43620 32866
rect 43740 32294 43860 32866
rect 44220 32294 44340 32866
rect 44474 32324 44596 32746
rect 44940 32340 45060 32760
rect 45404 32324 45526 32746
rect 45660 32294 45780 32866
rect 46140 32294 46260 32866
rect 46380 32310 46500 32730
rect 46620 32294 46740 32866
rect 46860 32294 46980 32866
rect 47670 32294 47790 32866
rect 48060 32294 48180 32866
rect 49110 32294 49230 32866
rect 49500 32294 49620 32866
rect 5340 31334 5460 31906
rect 5594 31454 5716 31876
rect 6060 31440 6180 31860
rect 6524 31454 6646 31876
rect 6780 31334 6900 31906
rect 7980 31334 8100 31906
rect 8220 31470 8340 31890
rect 8460 31334 8580 31906
rect 8700 31334 8820 31906
rect 9750 31334 9870 31906
rect 10140 31334 10260 31906
rect 11100 31334 11220 31906
rect 11354 31454 11476 31876
rect 11820 31440 11940 31860
rect 12284 31454 12406 31876
rect 12540 31334 12660 31906
rect 14700 31334 14820 31906
rect 14954 31454 15076 31876
rect 15420 31440 15540 31860
rect 15884 31454 16006 31876
rect 16140 31334 16260 31906
rect 17100 31334 17220 31906
rect 17354 31454 17476 31876
rect 17820 31440 17940 31860
rect 18284 31454 18406 31876
rect 18540 31334 18660 31906
rect 19260 31334 19380 31906
rect 19514 31454 19636 31876
rect 19980 31440 20100 31860
rect 20444 31454 20566 31876
rect 20700 31334 20820 31906
rect 21180 31334 21300 31906
rect 21570 31334 21690 31906
rect 22140 31334 22260 31906
rect 22380 31334 22500 31906
rect 22620 31470 22740 31890
rect 22860 31334 22980 31906
rect 23820 31650 23940 31920
rect 24060 31650 24180 31920
rect 24870 31634 24990 31906
rect 25110 31334 25230 31906
rect 25500 31334 25620 31906
rect 25980 31334 26100 31906
rect 26220 31334 26340 31906
rect 26460 31470 26580 31890
rect 26700 31334 26820 31906
rect 27180 31650 27300 31920
rect 27420 31650 27540 31920
rect 27750 31334 27870 31906
rect 28140 31334 28260 31906
rect 28620 31650 28740 31920
rect 28860 31650 28980 31920
rect 29100 31334 29220 31906
rect 29340 31334 29460 31906
rect 29580 31470 29700 31890
rect 29820 31334 29940 31906
rect 30780 31334 30900 31906
rect 31034 31454 31156 31876
rect 31500 31440 31620 31860
rect 31964 31454 32086 31876
rect 32220 31334 32340 31906
rect 33180 31334 33300 31906
rect 33570 31334 33690 31906
rect 34620 31334 34740 31906
rect 35010 31334 35130 31906
rect 36060 31334 36180 31906
rect 36300 31334 36420 31906
rect 36540 31470 36660 31890
rect 36780 31334 36900 31906
rect 37740 31334 37860 31906
rect 38130 31334 38250 31906
rect 38940 31334 39060 31906
rect 39180 31470 39300 31890
rect 39420 31334 39540 31906
rect 39660 31334 39780 31906
rect 40620 31650 40740 31920
rect 40860 31650 40980 31920
rect 41670 31334 41790 31906
rect 42060 31334 42180 31906
rect 43020 31334 43140 31906
rect 43260 31334 43380 31906
rect 43500 31470 43620 31890
rect 43740 31334 43860 31906
rect 44460 31334 44580 31906
rect 44700 31470 44820 31890
rect 44940 31334 45060 31906
rect 45180 31334 45300 31906
rect 46230 31334 46350 31906
rect 46620 31334 46740 31906
rect 48060 31334 48180 31906
rect 48314 31454 48436 31876
rect 48780 31440 48900 31860
rect 49244 31454 49366 31876
rect 49500 31334 49620 31906
rect 7020 26294 7140 26866
rect 7274 26324 7396 26746
rect 7740 26340 7860 26760
rect 8204 26324 8326 26746
rect 8460 26294 8580 26866
rect 8700 26294 8820 26866
rect 9090 26294 9210 26866
rect 9420 26294 9540 26866
rect 9674 26324 9796 26746
rect 10140 26340 10260 26760
rect 10604 26324 10726 26746
rect 10860 26294 10980 26866
rect 11100 26294 11220 26866
rect 11340 26310 11460 26730
rect 11580 26294 11700 26866
rect 11820 26294 11940 26866
rect 12060 26294 12180 26866
rect 12450 26294 12570 26866
rect 12780 26294 12900 26866
rect 13170 26294 13290 26866
rect 13830 26294 13950 26566
rect 14070 26294 14190 26866
rect 14460 26294 14580 26866
rect 15420 26294 15540 26866
rect 15810 26294 15930 26866
rect 16710 26294 16830 26866
rect 17100 26294 17220 26866
rect 18060 26294 18180 26866
rect 18450 26294 18570 26866
rect 19260 26294 19380 26866
rect 19500 26294 19620 26866
rect 19740 26310 19860 26730
rect 19980 26294 20100 26866
rect 20940 26294 21060 26866
rect 21330 26294 21450 26866
rect 22140 26294 22260 26866
rect 22530 26294 22650 26866
rect 23580 26294 23700 26866
rect 23970 26294 24090 26866
rect 25020 26294 25140 26866
rect 25410 26294 25530 26866
rect 26460 26294 26580 26866
rect 26850 26294 26970 26866
rect 28380 26294 28500 26866
rect 28620 26294 28740 26866
rect 28860 26310 28980 26730
rect 29100 26294 29220 26866
rect 30390 26294 30510 26866
rect 30780 26294 30900 26866
rect 31740 26294 31860 26866
rect 31980 26294 32100 26866
rect 32220 26310 32340 26730
rect 32460 26294 32580 26866
rect 32940 26294 33060 26866
rect 33194 26324 33316 26746
rect 33660 26340 33780 26760
rect 34124 26324 34246 26746
rect 34380 26294 34500 26866
rect 34860 26294 34980 26866
rect 35250 26294 35370 26866
rect 36060 26294 36180 26866
rect 36450 26294 36570 26866
rect 37590 26294 37710 26866
rect 37980 26294 38100 26866
rect 38700 26294 38820 26866
rect 39090 26294 39210 26866
rect 39660 26294 39780 26866
rect 39914 26324 40036 26746
rect 40380 26340 40500 26760
rect 40844 26324 40966 26746
rect 41100 26294 41220 26866
rect 41580 26294 41700 26866
rect 41970 26294 42090 26866
rect 43020 26294 43140 26866
rect 43260 26294 43380 26866
rect 43500 26310 43620 26730
rect 43740 26294 43860 26866
rect 44460 26294 44580 26866
rect 44700 26310 44820 26730
rect 44940 26294 45060 26866
rect 45180 26294 45300 26866
rect 45900 26294 46020 26866
rect 46140 26310 46260 26730
rect 46380 26294 46500 26866
rect 46620 26294 46740 26866
rect 46860 26280 46980 26550
rect 47100 26280 47220 26550
rect 47340 26294 47460 26866
rect 47790 26294 47910 26866
rect 48240 26294 48360 26866
rect 48540 26294 48660 26866
rect 48930 26294 49050 26866
rect 49260 26294 49380 26866
rect 49500 26310 49620 26730
rect 49740 26294 49860 26866
rect 49980 26294 50100 26866
rect 5340 25334 5460 25906
rect 5594 25454 5716 25876
rect 6060 25440 6180 25860
rect 6524 25454 6646 25876
rect 6780 25334 6900 25906
rect 7020 25334 7140 25906
rect 7410 25334 7530 25906
rect 7740 25334 7860 25906
rect 7980 25334 8100 25906
rect 8220 25470 8340 25890
rect 8460 25334 8580 25906
rect 8700 25334 8820 25906
rect 9090 25334 9210 25906
rect 9420 25334 9540 25906
rect 9674 25454 9796 25876
rect 10140 25440 10260 25860
rect 10604 25454 10726 25876
rect 10860 25334 10980 25906
rect 12060 25634 12180 25906
rect 12300 25334 12420 25906
rect 12690 25334 12810 25906
rect 13740 25650 13860 25920
rect 13980 25650 14100 25920
rect 14940 25334 15060 25906
rect 15180 25334 15300 25906
rect 15420 25470 15540 25890
rect 15660 25334 15780 25906
rect 20790 25334 20910 25906
rect 21180 25334 21300 25906
rect 23100 25334 23220 25906
rect 23490 25334 23610 25906
rect 25500 25334 25620 25906
rect 25754 25454 25876 25876
rect 26220 25440 26340 25860
rect 26684 25454 26806 25876
rect 26940 25334 27060 25906
rect 27900 25334 28020 25906
rect 28140 25334 28260 25906
rect 28380 25470 28500 25890
rect 28620 25334 28740 25906
rect 30300 25650 30420 25920
rect 30540 25650 30660 25920
rect 31020 25334 31140 25906
rect 31260 25334 31380 25906
rect 31500 25470 31620 25890
rect 31740 25334 31860 25906
rect 32220 25650 32340 25920
rect 32460 25650 32580 25920
rect 33180 25334 33300 25906
rect 33570 25334 33690 25906
rect 34620 25334 34740 25906
rect 35010 25334 35130 25906
rect 36060 25334 36180 25906
rect 36450 25334 36570 25906
rect 37500 25334 37620 25906
rect 37890 25334 38010 25906
rect 38940 25334 39060 25906
rect 39330 25334 39450 25906
rect 40380 25334 40500 25906
rect 40770 25334 40890 25906
rect 41820 25334 41940 25906
rect 42210 25334 42330 25906
rect 43260 25634 43380 25906
rect 43500 25634 43620 25906
rect 43740 25634 43860 25906
rect 44460 25650 44580 25920
rect 44700 25754 44820 25876
rect 47820 25334 47940 25906
rect 48074 25454 48196 25876
rect 48540 25440 48660 25860
rect 49004 25454 49126 25876
rect 49260 25334 49380 25906
rect 5340 20294 5460 20866
rect 5594 20324 5716 20746
rect 6060 20340 6180 20760
rect 6524 20324 6646 20746
rect 6780 20294 6900 20866
rect 8220 20294 8340 20866
rect 8610 20294 8730 20866
rect 9660 20294 9780 20866
rect 10050 20294 10170 20866
rect 11100 20294 11220 20866
rect 11340 20294 11460 20866
rect 11580 20310 11700 20730
rect 11820 20294 11940 20866
rect 14220 20294 14340 20866
rect 14474 20324 14596 20746
rect 14940 20340 15060 20760
rect 15404 20324 15526 20746
rect 15660 20294 15780 20866
rect 16860 20324 16980 20446
rect 17100 20280 17220 20550
rect 18060 20294 18180 20866
rect 18450 20294 18570 20866
rect 18780 20294 18900 20866
rect 19034 20324 19156 20746
rect 19500 20340 19620 20760
rect 19964 20324 20086 20746
rect 20220 20294 20340 20866
rect 20460 20294 20580 20866
rect 20714 20324 20836 20746
rect 21180 20340 21300 20760
rect 21644 20324 21766 20746
rect 21900 20294 22020 20866
rect 22140 20294 22260 20866
rect 22380 20294 22500 20866
rect 22620 20310 22740 20730
rect 22860 20294 22980 20866
rect 25020 20280 25140 20550
rect 25260 20280 25380 20550
rect 26220 20294 26340 20866
rect 26460 20294 26580 20866
rect 26700 20310 26820 20730
rect 26940 20294 27060 20866
rect 27900 20294 28020 20866
rect 28140 20294 28260 20866
rect 28380 20310 28500 20730
rect 28620 20294 28740 20866
rect 29100 20294 29220 20866
rect 29490 20294 29610 20866
rect 30300 20294 30420 20866
rect 30540 20310 30660 20730
rect 30780 20294 30900 20866
rect 31020 20294 31140 20866
rect 31980 20294 32100 20866
rect 32370 20294 32490 20866
rect 33180 20294 33300 20866
rect 33570 20294 33690 20866
rect 34620 20294 34740 20866
rect 35010 20294 35130 20866
rect 35820 20294 35940 20866
rect 36210 20294 36330 20866
rect 36780 20294 36900 20866
rect 37034 20324 37156 20746
rect 37500 20340 37620 20760
rect 37964 20324 38086 20746
rect 38220 20294 38340 20866
rect 38940 20294 39060 20866
rect 39180 20294 39300 20866
rect 39420 20310 39540 20730
rect 39660 20294 39780 20866
rect 40380 20294 40500 20866
rect 40770 20294 40890 20866
rect 41580 20294 41700 20866
rect 41820 20294 41940 20866
rect 42060 20310 42180 20730
rect 42300 20294 42420 20866
rect 43260 20294 43380 20566
rect 43500 20294 43620 20566
rect 43740 20294 43860 20566
rect 44220 20294 44340 20866
rect 44474 20324 44596 20746
rect 44940 20340 45060 20760
rect 45404 20324 45526 20746
rect 45660 20294 45780 20866
rect 45900 20294 46020 20866
rect 46154 20324 46276 20746
rect 46620 20340 46740 20760
rect 47084 20324 47206 20746
rect 47340 20294 47460 20866
rect 47580 20280 47700 20550
rect 47820 20280 47940 20550
rect 48780 20294 48900 20866
rect 49230 20294 49350 20866
rect 49680 20294 49800 20866
rect 5580 19334 5700 19906
rect 5820 19334 5940 19906
rect 6060 19470 6180 19890
rect 6300 19334 6420 19906
rect 8940 19334 9060 19906
rect 9194 19454 9316 19876
rect 9660 19440 9780 19860
rect 10124 19454 10246 19876
rect 10380 19334 10500 19906
rect 11580 19334 11700 19906
rect 11834 19454 11956 19876
rect 12300 19440 12420 19860
rect 12764 19454 12886 19876
rect 13020 19334 13140 19906
rect 13500 19334 13620 19906
rect 13754 19454 13876 19876
rect 14220 19440 14340 19860
rect 14684 19454 14806 19876
rect 14940 19334 15060 19906
rect 15510 19334 15630 19906
rect 15900 19334 16020 19906
rect 16140 19634 16260 19906
rect 17820 19334 17940 19906
rect 18060 19334 18180 19906
rect 18300 19470 18420 19890
rect 18540 19334 18660 19906
rect 19500 19334 19620 19906
rect 19890 19334 20010 19906
rect 20940 19334 21060 19906
rect 21330 19334 21450 19906
rect 22140 19334 22260 19906
rect 22530 19334 22650 19906
rect 23580 19334 23700 19906
rect 23970 19334 24090 19906
rect 24540 19334 24660 19906
rect 24794 19454 24916 19876
rect 25260 19440 25380 19860
rect 25724 19454 25846 19876
rect 25980 19334 26100 19906
rect 26220 19334 26340 19906
rect 26460 19470 26580 19890
rect 26700 19334 26820 19906
rect 26940 19334 27060 19906
rect 27180 19650 27300 19920
rect 27420 19650 27540 19920
rect 28380 19334 28500 19906
rect 28620 19334 28740 19906
rect 28860 19470 28980 19890
rect 29100 19334 29220 19906
rect 30540 19334 30660 19906
rect 30930 19334 31050 19906
rect 31980 19334 32100 19906
rect 32370 19334 32490 19906
rect 33180 19334 33300 19906
rect 33420 19470 33540 19890
rect 33660 19334 33780 19906
rect 33900 19334 34020 19906
rect 35820 19334 35940 19906
rect 36210 19334 36330 19906
rect 36780 19634 36900 19906
rect 37020 19334 37140 19906
rect 37410 19334 37530 19906
rect 37980 19334 38100 19906
rect 38370 19334 38490 19906
rect 38940 19334 39060 19906
rect 39330 19334 39450 19906
rect 40380 19334 40500 19906
rect 40770 19334 40890 19906
rect 41580 19650 41700 19920
rect 41820 19650 41940 19920
rect 42840 19334 42960 19906
rect 43290 19334 43410 19906
rect 43740 19334 43860 19906
rect 44460 19334 44580 19906
rect 44700 19470 44820 19890
rect 44940 19334 45060 19906
rect 45180 19334 45300 19906
rect 46140 19334 46260 19906
rect 46530 19334 46650 19906
rect 47580 19634 47700 19906
rect 47820 19634 47940 19906
rect 48060 19634 48180 19906
rect 49020 19334 49140 19906
rect 49260 19470 49380 19890
rect 49500 19334 49620 19906
rect 49740 19334 49860 19906
rect 6300 14294 6420 14866
rect 6690 14294 6810 14866
rect 7740 14294 7860 14866
rect 7994 14324 8116 14746
rect 8460 14340 8580 14760
rect 8924 14324 9046 14746
rect 9180 14294 9300 14866
rect 9420 14294 9540 14866
rect 9674 14324 9796 14746
rect 10140 14340 10260 14760
rect 10604 14324 10726 14746
rect 10860 14294 10980 14866
rect 11100 14294 11220 14866
rect 11354 14324 11476 14746
rect 11820 14340 11940 14760
rect 12284 14324 12406 14746
rect 12540 14294 12660 14866
rect 13260 14294 13380 14866
rect 13514 14324 13636 14746
rect 13980 14340 14100 14760
rect 14444 14324 14566 14746
rect 14700 14294 14820 14866
rect 14940 14294 15060 14866
rect 15194 14324 15316 14746
rect 15660 14340 15780 14760
rect 16124 14324 16246 14746
rect 16380 14294 16500 14866
rect 16710 14294 16830 14866
rect 17100 14294 17220 14866
rect 17340 14294 17460 14566
rect 17580 14280 17700 14550
rect 17820 14280 17940 14550
rect 18060 14294 18180 14866
rect 18300 14294 18420 14866
rect 18540 14310 18660 14730
rect 18780 14294 18900 14866
rect 19260 14294 19380 14866
rect 19650 14294 19770 14866
rect 20700 14294 20820 14866
rect 20940 14310 21060 14730
rect 21180 14294 21300 14866
rect 21420 14294 21540 14866
rect 22140 14294 22260 14866
rect 22380 14294 22500 14866
rect 22620 14310 22740 14730
rect 22860 14294 22980 14866
rect 23580 14294 23700 14866
rect 23970 14294 24090 14866
rect 24870 14294 24990 14866
rect 25260 14294 25380 14866
rect 25740 14294 25860 14866
rect 25994 14324 26116 14746
rect 26460 14340 26580 14760
rect 26924 14324 27046 14746
rect 27180 14294 27300 14866
rect 27900 14294 28020 14866
rect 28290 14294 28410 14866
rect 29100 14294 29220 14866
rect 29490 14294 29610 14866
rect 30300 14294 30420 14866
rect 30554 14324 30676 14746
rect 31020 14340 31140 14760
rect 31484 14324 31606 14746
rect 31740 14294 31860 14866
rect 32310 14294 32430 14866
rect 32700 14294 32820 14866
rect 33180 14294 33300 14866
rect 33570 14294 33690 14866
rect 34620 14294 34740 14866
rect 35010 14294 35130 14866
rect 36060 14294 36180 14866
rect 36300 14310 36420 14730
rect 36540 14294 36660 14866
rect 36780 14294 36900 14866
rect 37740 14294 37860 14866
rect 38130 14294 38250 14866
rect 38700 14294 38820 14866
rect 38954 14324 39076 14746
rect 39420 14340 39540 14760
rect 39884 14324 40006 14746
rect 40140 14294 40260 14866
rect 41580 14294 41700 14866
rect 41834 14324 41956 14746
rect 42300 14340 42420 14760
rect 42764 14324 42886 14746
rect 43020 14294 43140 14866
rect 44460 14294 44580 14866
rect 44700 14310 44820 14730
rect 44940 14294 45060 14866
rect 45180 14294 45300 14866
rect 46140 14294 46260 14866
rect 46530 14294 46650 14866
rect 47670 14294 47790 14866
rect 48060 14294 48180 14866
rect 49020 14294 49140 14866
rect 49260 14310 49380 14730
rect 49500 14294 49620 14866
rect 49740 14294 49860 14866
rect 6870 13334 6990 13906
rect 7260 13334 7380 13906
rect 8940 13334 9060 13906
rect 9180 13470 9300 13890
rect 9420 13334 9540 13906
rect 9660 13320 9780 13740
rect 9900 13334 10020 13906
rect 10860 13334 10980 13906
rect 11250 13334 11370 13906
rect 12060 13334 12180 13906
rect 12300 13334 12420 13906
rect 12540 13470 12660 13890
rect 12780 13334 12900 13906
rect 15900 13334 16020 13906
rect 16290 13334 16410 13906
rect 16620 13334 16740 13906
rect 16860 13334 16980 13906
rect 17100 13470 17220 13890
rect 17340 13334 17460 13906
rect 17580 13334 17700 13906
rect 17834 13454 17956 13876
rect 18300 13440 18420 13860
rect 18764 13454 18886 13876
rect 19020 13334 19140 13906
rect 19260 13334 19380 13906
rect 19514 13454 19636 13876
rect 19980 13440 20100 13860
rect 20444 13454 20566 13876
rect 20700 13334 20820 13906
rect 21900 13334 22020 13906
rect 22154 13454 22276 13876
rect 22620 13440 22740 13860
rect 23084 13454 23206 13876
rect 23340 13334 23460 13906
rect 25020 13334 25140 13906
rect 25260 13470 25380 13890
rect 25500 13334 25620 13906
rect 25740 13334 25860 13906
rect 26700 13334 26820 13906
rect 27090 13334 27210 13906
rect 29100 13334 29220 13906
rect 29340 13470 29460 13890
rect 29580 13334 29700 13906
rect 29820 13334 29940 13906
rect 30300 13334 30420 13906
rect 30540 13334 30660 13906
rect 30780 13470 30900 13890
rect 31020 13334 31140 13906
rect 32070 13334 32190 13906
rect 32460 13334 32580 13906
rect 32940 13334 33060 13906
rect 33194 13454 33316 13876
rect 33660 13440 33780 13860
rect 34124 13454 34246 13876
rect 34380 13334 34500 13906
rect 34620 13334 34740 13906
rect 34860 13470 34980 13890
rect 35100 13334 35220 13906
rect 35340 13334 35460 13906
rect 36060 13334 36180 13906
rect 36450 13334 36570 13906
rect 37500 13334 37620 13906
rect 37890 13334 38010 13906
rect 38940 13334 39060 13906
rect 39330 13334 39450 13906
rect 40140 13334 40260 13906
rect 40380 13334 40500 13906
rect 40620 13470 40740 13890
rect 40860 13334 40980 13906
rect 41580 13334 41700 13906
rect 41970 13334 42090 13906
rect 42210 13634 42330 13906
rect 43260 13334 43380 13906
rect 43650 13334 43770 13906
rect 44460 13334 44580 13906
rect 44700 13470 44820 13890
rect 44940 13334 45060 13906
rect 45180 13334 45300 13906
rect 46140 13334 46260 13906
rect 46530 13334 46650 13906
rect 47580 13334 47700 13906
rect 47820 13470 47940 13890
rect 48060 13334 48180 13906
rect 48300 13334 48420 13906
rect 49350 13334 49470 13906
rect 49740 13334 49860 13906
rect 5580 8294 5700 8866
rect 5820 8294 5940 8866
rect 6060 8310 6180 8730
rect 6300 8294 6420 8866
rect 6780 8294 6900 8866
rect 7170 8294 7290 8866
rect 7740 8294 7860 8866
rect 7994 8324 8116 8746
rect 8460 8340 8580 8760
rect 8924 8324 9046 8746
rect 9180 8294 9300 8866
rect 9750 8294 9870 8566
rect 9990 8294 10110 8866
rect 10380 8294 10500 8866
rect 11430 8294 11550 8866
rect 11820 8294 11940 8866
rect 13740 8294 13860 8866
rect 13994 8324 14116 8746
rect 14460 8340 14580 8760
rect 14924 8324 15046 8746
rect 15180 8294 15300 8866
rect 16380 8294 16500 8866
rect 16770 8294 16890 8866
rect 17340 8294 17460 8866
rect 17594 8324 17716 8746
rect 18060 8340 18180 8760
rect 18524 8324 18646 8746
rect 18780 8294 18900 8866
rect 19260 8294 19380 8866
rect 19514 8324 19636 8746
rect 19980 8340 20100 8760
rect 20444 8324 20566 8746
rect 20700 8294 20820 8866
rect 21270 8294 21390 8866
rect 21660 8294 21780 8866
rect 21900 8294 22020 8866
rect 22154 8324 22276 8746
rect 22620 8340 22740 8760
rect 23084 8324 23206 8746
rect 23340 8294 23460 8866
rect 23820 8294 23940 8866
rect 24210 8294 24330 8866
rect 25500 8294 25620 8866
rect 25754 8324 25876 8746
rect 26220 8340 26340 8760
rect 26684 8324 26806 8746
rect 26940 8294 27060 8866
rect 27900 8294 28020 8866
rect 28290 8294 28410 8866
rect 29340 8280 29460 8550
rect 29580 8280 29700 8550
rect 30540 8280 30660 8550
rect 30780 8280 30900 8550
rect 31740 8294 31860 8866
rect 31980 8310 32100 8730
rect 32220 8294 32340 8866
rect 32460 8294 32580 8866
rect 33180 8294 33300 8866
rect 33434 8324 33556 8746
rect 33900 8340 34020 8760
rect 34364 8324 34486 8746
rect 34620 8294 34740 8866
rect 35670 8294 35790 8566
rect 35910 8294 36030 8866
rect 36300 8294 36420 8866
rect 36780 8294 36900 8866
rect 37170 8294 37290 8866
rect 37830 8294 37950 8566
rect 38070 8294 38190 8866
rect 38460 8294 38580 8866
rect 38940 8294 39060 8866
rect 39180 8310 39300 8730
rect 39420 8294 39540 8866
rect 39660 8294 39780 8866
rect 40380 8294 40500 8866
rect 40770 8294 40890 8866
rect 41580 8294 41700 8866
rect 41970 8294 42090 8866
rect 42540 8294 42660 8866
rect 42794 8324 42916 8746
rect 43260 8340 43380 8760
rect 43724 8324 43846 8746
rect 43980 8294 44100 8866
rect 45180 8294 45300 8866
rect 45434 8324 45556 8746
rect 45900 8340 46020 8760
rect 46364 8324 46486 8746
rect 46620 8294 46740 8866
rect 47670 8294 47790 8866
rect 48060 8294 48180 8866
rect 49110 8294 49230 8866
rect 49500 8294 49620 8866
rect 5580 7334 5700 7906
rect 5834 7454 5956 7876
rect 6300 7440 6420 7860
rect 6764 7454 6886 7876
rect 7020 7334 7140 7906
rect 7980 7650 8100 7920
rect 8220 7650 8340 7920
rect 8700 7334 8820 7906
rect 8940 7334 9060 7906
rect 9180 7470 9300 7890
rect 9420 7334 9540 7906
rect 9900 7334 10020 7906
rect 10290 7334 10410 7906
rect 10860 7334 10980 7906
rect 11100 7334 11220 7906
rect 11340 7470 11460 7890
rect 11580 7334 11700 7906
rect 12300 7334 12420 7906
rect 12690 7334 12810 7906
rect 13830 7334 13950 7906
rect 14220 7334 14340 7906
rect 14460 7634 14580 7906
rect 15420 7634 15540 7906
rect 15660 7634 15780 7906
rect 15900 7634 16020 7906
rect 18060 7634 18180 7906
rect 18300 7634 18420 7906
rect 18540 7634 18660 7906
rect 20700 7334 20820 7906
rect 21090 7334 21210 7906
rect 23340 7334 23460 7906
rect 23730 7334 23850 7906
rect 25740 7334 25860 7906
rect 25994 7454 26116 7876
rect 26460 7440 26580 7860
rect 26924 7454 27046 7876
rect 27180 7334 27300 7906
rect 27900 7334 28020 7906
rect 28290 7334 28410 7906
rect 29100 7334 29220 7906
rect 29490 7334 29610 7906
rect 30060 7334 30180 7906
rect 30314 7454 30436 7876
rect 30780 7440 30900 7860
rect 31244 7454 31366 7876
rect 31500 7334 31620 7906
rect 31980 7334 32100 7906
rect 32220 7470 32340 7890
rect 32460 7334 32580 7906
rect 32700 7334 32820 7906
rect 33180 7334 33300 7906
rect 33570 7334 33690 7906
rect 34710 7334 34830 7906
rect 35100 7334 35220 7906
rect 36060 7334 36180 7906
rect 36450 7334 36570 7906
rect 37500 7334 37620 7906
rect 37740 7334 37860 7906
rect 37980 7470 38100 7890
rect 38220 7334 38340 7906
rect 38940 7334 39060 7906
rect 39330 7334 39450 7906
rect 40380 7334 40500 7906
rect 40770 7334 40890 7906
rect 43260 7634 43380 7906
rect 43500 7634 43620 7906
rect 43740 7634 43860 7906
rect 44520 7334 44640 7906
rect 44970 7334 45090 7906
rect 45420 7334 45540 7906
rect 46380 7650 46500 7920
rect 46620 7650 46740 7920
rect 47340 7334 47460 7906
rect 47580 7334 47700 7906
rect 47820 7470 47940 7890
rect 48060 7334 48180 7906
<< pdcontact >>
rect 5670 41294 5790 41866
rect 5910 41294 6030 42466
rect 6300 41294 6420 42466
rect 6780 41294 6900 41866
rect 7020 41294 7140 41866
rect 7260 41294 7380 41866
rect 7830 41294 7950 41866
rect 8070 41294 8190 42466
rect 8460 41294 8580 42466
rect 8940 41294 9060 42466
rect 9194 41340 9316 42210
rect 9660 41294 9780 42466
rect 10124 41340 10246 42210
rect 10380 41294 10500 42466
rect 10950 41310 11070 42480
rect 11340 41310 11460 42480
rect 12390 41310 12510 42480
rect 12780 41310 12900 42480
rect 13740 41294 13860 42466
rect 14130 41294 14250 42466
rect 14370 41294 14490 41866
rect 15420 41294 15540 41866
rect 15660 41294 15780 41866
rect 15900 41294 16020 41866
rect 17100 41294 17220 42466
rect 17490 41294 17610 42466
rect 17730 41294 17850 41866
rect 19260 41294 19380 42466
rect 19514 41340 19636 42210
rect 19980 41294 20100 42466
rect 20444 41340 20566 42210
rect 20700 41294 20820 42466
rect 21180 41310 21300 41880
rect 21420 41310 21540 41880
rect 22620 41294 22740 42466
rect 22874 41340 22996 42210
rect 23340 41294 23460 42466
rect 23804 41340 23926 42210
rect 24060 41294 24180 42466
rect 25110 41294 25230 41866
rect 25350 41294 25470 42466
rect 25740 41294 25860 42466
rect 26700 41294 26820 41866
rect 26940 41294 27060 41866
rect 27180 41294 27300 41866
rect 27900 41294 28020 42466
rect 28290 41294 28410 42466
rect 28530 41294 28650 41866
rect 29100 41294 29220 41866
rect 29340 41294 29460 41866
rect 29580 41294 29700 41866
rect 30300 41294 30420 42466
rect 30690 41294 30810 42466
rect 30930 41294 31050 41866
rect 31740 41294 31860 42466
rect 32130 41294 32250 42466
rect 32370 41294 32490 41866
rect 33180 41294 33300 41866
rect 33420 41294 33540 41866
rect 33660 41294 33780 41866
rect 34620 41310 34740 42480
rect 35010 41310 35130 42480
rect 35820 41294 35940 42466
rect 36074 41340 36196 42210
rect 36540 41294 36660 42466
rect 37004 41340 37126 42210
rect 37260 41294 37380 42466
rect 37830 41294 37950 41866
rect 38070 41294 38190 42466
rect 38460 41294 38580 42466
rect 39420 41294 39540 42466
rect 39674 41340 39796 42210
rect 40140 41294 40260 42466
rect 40604 41340 40726 42210
rect 40860 41294 40980 42466
rect 41820 41310 41940 41880
rect 42060 41310 42180 41880
rect 43020 41294 43140 42466
rect 43410 41294 43530 42466
rect 43650 41294 43770 41866
rect 44220 41294 44340 42466
rect 44610 41294 44730 42466
rect 44850 41294 44970 41866
rect 45180 41310 45300 41880
rect 45420 41310 45540 41880
rect 45660 41294 45780 42466
rect 45914 41340 46036 42210
rect 46380 41294 46500 42466
rect 46844 41340 46966 42210
rect 47100 41294 47220 42466
rect 47340 41294 47460 42466
rect 47594 41340 47716 42210
rect 48060 41294 48180 42466
rect 48524 41340 48646 42210
rect 48780 41294 48900 42466
rect 5820 39854 5940 40876
rect 6060 39900 6180 40920
rect 6300 39734 6420 40906
rect 6540 39734 6660 40906
rect 8220 40334 8340 40906
rect 8460 40334 8580 40906
rect 8700 40334 8820 40906
rect 9660 40334 9780 40906
rect 9900 40334 10020 40906
rect 10140 40334 10260 40906
rect 10620 39734 10740 40906
rect 10860 39734 10980 40906
rect 11100 39900 11220 40920
rect 11340 39854 11460 40876
rect 11580 39734 11700 40906
rect 11834 39990 11956 40860
rect 12300 39734 12420 40906
rect 12764 39990 12886 40860
rect 13020 39734 13140 40906
rect 13500 40334 13620 40906
rect 13740 40334 13860 40906
rect 13980 40334 14100 40906
rect 14460 40334 14580 40906
rect 14700 40334 14820 40906
rect 14940 40334 15060 40906
rect 15180 40334 15300 40906
rect 15660 40320 15780 40890
rect 15900 40320 16020 40890
rect 16380 39734 16500 40906
rect 16770 39734 16890 40906
rect 17010 40334 17130 40906
rect 17670 40334 17790 40906
rect 17910 39734 18030 40906
rect 18300 39734 18420 40906
rect 18540 40320 18660 40890
rect 18780 40320 18900 40890
rect 19260 39734 19380 40906
rect 19650 39734 19770 40906
rect 19890 40334 20010 40906
rect 20940 40334 21060 40906
rect 21180 40334 21300 40906
rect 21420 40334 21540 40906
rect 21900 39734 22020 40906
rect 22154 39990 22276 40860
rect 22620 39734 22740 40906
rect 23084 39990 23206 40860
rect 23340 39734 23460 40906
rect 23820 39720 23940 40890
rect 24210 39720 24330 40890
rect 24780 39734 24900 40906
rect 25170 39734 25290 40906
rect 25410 40334 25530 40906
rect 26220 39854 26340 40876
rect 26460 39900 26580 40920
rect 26700 39734 26820 40906
rect 26940 39720 27060 40740
rect 27180 39734 27300 40906
rect 27900 40320 28020 40890
rect 28140 40320 28260 40890
rect 30540 40334 30660 40906
rect 30780 40334 30900 40906
rect 31020 40334 31140 40906
rect 31980 40334 32100 40906
rect 32220 40334 32340 40906
rect 32460 40334 32580 40906
rect 33420 39734 33540 40906
rect 33674 39990 33796 40860
rect 34140 39734 34260 40906
rect 34604 39990 34726 40860
rect 34860 39734 34980 40906
rect 36060 39734 36180 40906
rect 36450 39734 36570 40906
rect 36690 40334 36810 40906
rect 37740 40334 37860 40906
rect 37980 40334 38100 40906
rect 38220 40334 38340 40906
rect 38940 39734 39060 40906
rect 39330 39734 39450 40906
rect 39570 40334 39690 40906
rect 40380 40334 40500 40906
rect 40620 40334 40740 40906
rect 40860 40334 40980 40906
rect 41820 40320 41940 40890
rect 42060 40320 42180 40890
rect 43020 39734 43140 40906
rect 43410 39734 43530 40906
rect 43650 40334 43770 40906
rect 44700 40320 44820 40890
rect 44940 40320 45060 40890
rect 45990 40334 46110 40906
rect 46230 39734 46350 40906
rect 46620 39734 46740 40906
rect 47580 39734 47700 40906
rect 47970 39734 48090 40906
rect 48210 40334 48330 40906
rect 49260 40334 49380 40906
rect 49500 40334 49620 40906
rect 49740 40334 49860 40906
rect 5580 35294 5700 35866
rect 5820 35294 5940 35866
rect 6060 35294 6180 35866
rect 7020 35310 7140 35880
rect 7260 35310 7380 35880
rect 8310 35294 8430 35866
rect 8550 35294 8670 36466
rect 8940 35294 9060 36466
rect 10860 35294 10980 35866
rect 11100 35294 11220 35866
rect 11340 35294 11460 35866
rect 12150 35294 12270 35866
rect 12390 35294 12510 36466
rect 12780 35294 12900 36466
rect 15030 35294 15150 35866
rect 15270 35294 15390 36466
rect 15660 35294 15780 36466
rect 16620 35294 16740 35866
rect 16860 35294 16980 35866
rect 17100 35294 17220 35866
rect 17340 35294 17460 35866
rect 18060 35294 18180 35866
rect 18300 35294 18420 35866
rect 18540 35294 18660 35866
rect 19500 35294 19620 35866
rect 19740 35294 19860 35866
rect 19980 35294 20100 35866
rect 20940 35294 21060 35866
rect 21180 35294 21300 35866
rect 21420 35294 21540 35866
rect 22380 35294 22500 35866
rect 22620 35294 22740 35866
rect 22860 35294 22980 35866
rect 23820 35310 23940 35880
rect 24060 35310 24180 35880
rect 25020 35294 25140 35866
rect 25260 35294 25380 35866
rect 25500 35294 25620 35866
rect 26460 35294 26580 36466
rect 26850 35294 26970 36466
rect 27090 35294 27210 35866
rect 27900 35294 28020 35866
rect 28140 35294 28260 35866
rect 28380 35294 28500 35866
rect 29100 35294 29220 35866
rect 29340 35294 29460 35866
rect 29580 35294 29700 35866
rect 30060 35294 30180 36466
rect 30450 35294 30570 36466
rect 30690 35294 30810 35866
rect 31260 35310 31380 35880
rect 31500 35310 31620 35880
rect 32070 35294 32190 35866
rect 32310 35294 32430 36466
rect 32700 35294 32820 36466
rect 33180 35294 33300 35866
rect 33420 35294 33540 35866
rect 33660 35294 33780 35866
rect 34620 35294 34740 35866
rect 34860 35294 34980 35866
rect 35100 35294 35220 35866
rect 35580 35294 35700 36466
rect 35834 35340 35956 36210
rect 36300 35294 36420 36466
rect 36764 35340 36886 36210
rect 37020 35294 37140 36466
rect 38940 35310 39060 35880
rect 39180 35310 39300 35880
rect 39900 35294 40020 36466
rect 40140 35460 40260 36480
rect 40380 35294 40500 36466
rect 40620 35280 40740 36300
rect 40860 35324 40980 36346
rect 41580 35310 41700 35880
rect 41820 35310 41940 35880
rect 42390 35294 42510 35866
rect 42630 35294 42750 36466
rect 43020 35294 43140 36466
rect 43500 35310 43620 35880
rect 43740 35310 43860 35880
rect 44460 35294 44580 36466
rect 44850 35294 44970 36466
rect 45090 35294 45210 35866
rect 46140 35294 46260 35866
rect 46380 35294 46500 35866
rect 46620 35294 46740 35866
rect 47580 35294 47700 36466
rect 47970 35294 48090 36466
rect 48210 35294 48330 35866
rect 49260 35294 49380 35866
rect 49500 35294 49620 35866
rect 49740 35294 49860 35866
rect 6630 34334 6750 34906
rect 6870 33734 6990 34906
rect 7260 33734 7380 34906
rect 7830 34334 7950 34906
rect 8070 33734 8190 34906
rect 8460 33734 8580 34906
rect 8940 33734 9060 34906
rect 9194 33990 9316 34860
rect 9660 33734 9780 34906
rect 10124 33990 10246 34860
rect 10380 33734 10500 34906
rect 11100 33734 11220 34906
rect 11354 33990 11476 34860
rect 11820 33734 11940 34906
rect 12284 33990 12406 34860
rect 12540 33734 12660 34906
rect 13740 34320 13860 34890
rect 13980 34320 14100 34890
rect 15180 34334 15300 34906
rect 15420 34334 15540 34906
rect 15660 34334 15780 34906
rect 16620 33734 16740 34906
rect 17010 33734 17130 34906
rect 17250 34334 17370 34906
rect 19260 34334 19380 34906
rect 19500 34334 19620 34906
rect 19740 34334 19860 34906
rect 20700 34334 20820 34906
rect 20940 34334 21060 34906
rect 21180 34334 21300 34906
rect 21420 34334 21540 34906
rect 23340 33734 23460 34906
rect 23730 33734 23850 34906
rect 23970 34334 24090 34906
rect 24780 33734 24900 34906
rect 25170 33734 25290 34906
rect 25410 34334 25530 34906
rect 25980 33734 26100 34906
rect 26234 33990 26356 34860
rect 26700 33734 26820 34906
rect 27164 33990 27286 34860
rect 27420 33734 27540 34906
rect 30300 34320 30420 34890
rect 30540 34320 30660 34890
rect 31020 34334 31140 34906
rect 31260 34334 31380 34906
rect 31500 34334 31620 34906
rect 31980 33734 32100 34906
rect 32370 33734 32490 34906
rect 32610 34334 32730 34906
rect 33180 34334 33300 34906
rect 33420 34334 33540 34906
rect 33660 34334 33780 34906
rect 34620 34334 34740 34906
rect 34860 34334 34980 34906
rect 35100 34334 35220 34906
rect 36060 34334 36180 34906
rect 36300 34334 36420 34906
rect 36540 34334 36660 34906
rect 37500 34334 37620 34906
rect 37740 34334 37860 34906
rect 37980 34334 38100 34906
rect 38940 34334 39060 34906
rect 39180 34334 39300 34906
rect 39420 34334 39540 34906
rect 40140 33734 40260 34906
rect 40530 33734 40650 34906
rect 40770 34334 40890 34906
rect 41580 34334 41700 34906
rect 41820 34334 41940 34906
rect 42060 34334 42180 34906
rect 43020 33734 43140 34906
rect 43410 33734 43530 34906
rect 43650 34334 43770 34906
rect 44220 33734 44340 34906
rect 44474 33990 44596 34860
rect 44940 33734 45060 34906
rect 45404 33990 45526 34860
rect 45660 33734 45780 34906
rect 46140 33734 46260 34906
rect 46530 33734 46650 34906
rect 46770 34334 46890 34906
rect 47580 34334 47700 34906
rect 47820 34334 47940 34906
rect 48060 34334 48180 34906
rect 49020 34334 49140 34906
rect 49260 34334 49380 34906
rect 49500 34334 49620 34906
rect 5340 29294 5460 30466
rect 5594 29340 5716 30210
rect 6060 29294 6180 30466
rect 6524 29340 6646 30210
rect 6780 29294 6900 30466
rect 7980 29294 8100 30466
rect 8370 29294 8490 30466
rect 8610 29294 8730 29866
rect 9660 29294 9780 29866
rect 9900 29294 10020 29866
rect 10140 29294 10260 29866
rect 11100 29294 11220 30466
rect 11354 29340 11476 30210
rect 11820 29294 11940 30466
rect 12284 29340 12406 30210
rect 12540 29294 12660 30466
rect 14700 29294 14820 30466
rect 14954 29340 15076 30210
rect 15420 29294 15540 30466
rect 15884 29340 16006 30210
rect 16140 29294 16260 30466
rect 17100 29294 17220 30466
rect 17354 29340 17476 30210
rect 17820 29294 17940 30466
rect 18284 29340 18406 30210
rect 18540 29294 18660 30466
rect 19260 29294 19380 30466
rect 19514 29340 19636 30210
rect 19980 29294 20100 30466
rect 20444 29340 20566 30210
rect 20700 29294 20820 30466
rect 21180 29294 21300 29866
rect 21420 29294 21540 29866
rect 21660 29294 21780 29866
rect 22230 29294 22350 29866
rect 22470 29294 22590 30466
rect 22860 29294 22980 30466
rect 23820 29310 23940 29880
rect 24060 29310 24180 29880
rect 24780 29294 24900 29866
rect 25020 29294 25140 29866
rect 25260 29294 25380 29866
rect 25500 29294 25620 29866
rect 26070 29294 26190 29866
rect 26310 29294 26430 30466
rect 26700 29294 26820 30466
rect 27180 29310 27300 29880
rect 27420 29310 27540 29880
rect 27660 29294 27780 29866
rect 27900 29294 28020 29866
rect 28140 29294 28260 29866
rect 28620 29310 28740 29880
rect 28860 29310 28980 29880
rect 29190 29294 29310 29866
rect 29430 29294 29550 30466
rect 29820 29294 29940 30466
rect 30780 29294 30900 30466
rect 31034 29340 31156 30210
rect 31500 29294 31620 30466
rect 31964 29340 32086 30210
rect 32220 29294 32340 30466
rect 33180 29294 33300 29866
rect 33420 29294 33540 29866
rect 33660 29294 33780 29866
rect 34620 29294 34740 29866
rect 34860 29294 34980 29866
rect 35100 29294 35220 29866
rect 36150 29294 36270 29866
rect 36390 29294 36510 30466
rect 36780 29294 36900 30466
rect 37740 29294 37860 29866
rect 37980 29294 38100 29866
rect 38220 29294 38340 29866
rect 38940 29294 39060 30466
rect 39330 29294 39450 30466
rect 39570 29294 39690 29866
rect 40620 29310 40740 29880
rect 40860 29310 40980 29880
rect 41580 29294 41700 29866
rect 41820 29294 41940 29866
rect 42060 29294 42180 29866
rect 43110 29294 43230 29866
rect 43350 29294 43470 30466
rect 43740 29294 43860 30466
rect 44460 29294 44580 30466
rect 44850 29294 44970 30466
rect 45090 29294 45210 29866
rect 46140 29294 46260 29866
rect 46380 29294 46500 29866
rect 46620 29294 46740 29866
rect 48060 29294 48180 30466
rect 48314 29340 48436 30210
rect 48780 29294 48900 30466
rect 49244 29340 49366 30210
rect 49500 29294 49620 30466
rect 7020 27734 7140 28906
rect 7274 27990 7396 28860
rect 7740 27734 7860 28906
rect 8204 27990 8326 28860
rect 8460 27734 8580 28906
rect 8700 28334 8820 28906
rect 8940 28334 9060 28906
rect 9180 28334 9300 28906
rect 9420 27734 9540 28906
rect 9674 27990 9796 28860
rect 10140 27734 10260 28906
rect 10604 27990 10726 28860
rect 10860 27734 10980 28906
rect 11100 27734 11220 28906
rect 11490 27734 11610 28906
rect 11730 28334 11850 28906
rect 12060 28334 12180 28906
rect 12300 28334 12420 28906
rect 12540 28334 12660 28906
rect 12780 28334 12900 28906
rect 13020 28334 13140 28906
rect 13260 28334 13380 28906
rect 13740 28334 13860 28906
rect 13980 28334 14100 28906
rect 14220 28334 14340 28906
rect 14460 28334 14580 28906
rect 15420 28334 15540 28906
rect 15660 28334 15780 28906
rect 15900 28334 16020 28906
rect 16620 28334 16740 28906
rect 16860 28334 16980 28906
rect 17100 28334 17220 28906
rect 18060 28334 18180 28906
rect 18300 28334 18420 28906
rect 18540 28334 18660 28906
rect 19350 28334 19470 28906
rect 19590 27734 19710 28906
rect 19980 27734 20100 28906
rect 20940 28334 21060 28906
rect 21180 28334 21300 28906
rect 21420 28334 21540 28906
rect 22140 28334 22260 28906
rect 22380 28334 22500 28906
rect 22620 28334 22740 28906
rect 23580 28334 23700 28906
rect 23820 28334 23940 28906
rect 24060 28334 24180 28906
rect 25020 28334 25140 28906
rect 25260 28334 25380 28906
rect 25500 28334 25620 28906
rect 26460 28334 26580 28906
rect 26700 28334 26820 28906
rect 26940 28334 27060 28906
rect 28470 28334 28590 28906
rect 28710 27734 28830 28906
rect 29100 27734 29220 28906
rect 30300 28334 30420 28906
rect 30540 28334 30660 28906
rect 30780 28334 30900 28906
rect 31830 28334 31950 28906
rect 32070 27734 32190 28906
rect 32460 27734 32580 28906
rect 32940 27734 33060 28906
rect 33194 27990 33316 28860
rect 33660 27734 33780 28906
rect 34124 27990 34246 28860
rect 34380 27734 34500 28906
rect 34860 28334 34980 28906
rect 35100 28334 35220 28906
rect 35340 28334 35460 28906
rect 36060 28334 36180 28906
rect 36300 28334 36420 28906
rect 36540 28334 36660 28906
rect 37500 28334 37620 28906
rect 37740 28334 37860 28906
rect 37980 28334 38100 28906
rect 38700 28334 38820 28906
rect 38940 28334 39060 28906
rect 39180 28334 39300 28906
rect 39660 27734 39780 28906
rect 39914 27990 40036 28860
rect 40380 27734 40500 28906
rect 40844 27990 40966 28860
rect 41100 27734 41220 28906
rect 41580 28334 41700 28906
rect 41820 28334 41940 28906
rect 42060 28334 42180 28906
rect 43110 28334 43230 28906
rect 43350 27734 43470 28906
rect 43740 27734 43860 28906
rect 44460 27734 44580 28906
rect 44850 27734 44970 28906
rect 45090 28334 45210 28906
rect 45900 27734 46020 28906
rect 46290 27734 46410 28906
rect 46530 28334 46650 28906
rect 46860 28320 46980 28890
rect 47100 28320 47220 28890
rect 47340 27734 47460 28906
rect 47580 27720 47700 28740
rect 47820 27734 47940 28906
rect 48060 27900 48180 28920
rect 48300 27854 48420 28876
rect 48540 28334 48660 28906
rect 48780 28334 48900 28906
rect 49020 28334 49140 28906
rect 49260 27734 49380 28906
rect 49650 27734 49770 28906
rect 49890 28334 50010 28906
rect 5340 23294 5460 24466
rect 5594 23340 5716 24210
rect 6060 23294 6180 24466
rect 6524 23340 6646 24210
rect 6780 23294 6900 24466
rect 7020 23294 7140 23866
rect 7260 23294 7380 23866
rect 7500 23294 7620 23866
rect 7830 23294 7950 23866
rect 8070 23294 8190 24466
rect 8460 23294 8580 24466
rect 8700 23294 8820 23866
rect 8940 23294 9060 23866
rect 9180 23294 9300 23866
rect 9420 23294 9540 24466
rect 9674 23340 9796 24210
rect 10140 23294 10260 24466
rect 10604 23340 10726 24210
rect 10860 23294 10980 24466
rect 12060 23294 12180 24466
rect 12300 23294 12420 24466
rect 12540 23280 12660 24300
rect 12780 23324 12900 24346
rect 13740 23310 13860 23880
rect 13980 23310 14100 23880
rect 15030 23294 15150 23866
rect 15270 23294 15390 24466
rect 15660 23294 15780 24466
rect 20700 23294 20820 23866
rect 20940 23294 21060 23866
rect 21180 23294 21300 23866
rect 23100 23294 23220 23866
rect 23340 23294 23460 23866
rect 23580 23294 23700 23866
rect 25500 23294 25620 24466
rect 25754 23340 25876 24210
rect 26220 23294 26340 24466
rect 26684 23340 26806 24210
rect 26940 23294 27060 24466
rect 27990 23294 28110 23866
rect 28230 23294 28350 24466
rect 28620 23294 28740 24466
rect 30300 23310 30420 23880
rect 30540 23310 30660 23880
rect 31110 23294 31230 23866
rect 31350 23294 31470 24466
rect 31740 23294 31860 24466
rect 32220 23310 32340 23880
rect 32460 23310 32580 23880
rect 33180 23294 33300 23866
rect 33420 23294 33540 23866
rect 33660 23294 33780 23866
rect 34620 23294 34740 23866
rect 34860 23294 34980 23866
rect 35100 23294 35220 23866
rect 36060 23294 36180 23866
rect 36300 23294 36420 23866
rect 36540 23294 36660 23866
rect 37500 23294 37620 23866
rect 37740 23294 37860 23866
rect 37980 23294 38100 23866
rect 38940 23294 39060 23866
rect 39180 23294 39300 23866
rect 39420 23294 39540 23866
rect 40380 23294 40500 23866
rect 40620 23294 40740 23866
rect 40860 23294 40980 23866
rect 41820 23294 41940 23866
rect 42060 23294 42180 23866
rect 42300 23294 42420 23866
rect 43260 23310 43380 24480
rect 43650 23310 43770 24480
rect 44460 23310 44580 23880
rect 44700 23310 44820 23880
rect 47820 23294 47940 24466
rect 48074 23340 48196 24210
rect 48540 23294 48660 24466
rect 49004 23340 49126 24210
rect 49260 23294 49380 24466
rect 5340 21734 5460 22906
rect 5594 21990 5716 22860
rect 6060 21734 6180 22906
rect 6524 21990 6646 22860
rect 6780 21734 6900 22906
rect 8220 22334 8340 22906
rect 8460 22334 8580 22906
rect 8700 22334 8820 22906
rect 9660 22334 9780 22906
rect 9900 22334 10020 22906
rect 10140 22334 10260 22906
rect 11190 22334 11310 22906
rect 11430 21734 11550 22906
rect 11820 21734 11940 22906
rect 14220 21734 14340 22906
rect 14474 21990 14596 22860
rect 14940 21734 15060 22906
rect 15404 21990 15526 22860
rect 15660 21734 15780 22906
rect 16860 22320 16980 22890
rect 17100 22320 17220 22890
rect 18060 22334 18180 22906
rect 18300 22334 18420 22906
rect 18540 22334 18660 22906
rect 18780 21734 18900 22906
rect 19034 21990 19156 22860
rect 19500 21734 19620 22906
rect 19964 21990 20086 22860
rect 20220 21734 20340 22906
rect 20460 21734 20580 22906
rect 20714 21990 20836 22860
rect 21180 21734 21300 22906
rect 21644 21990 21766 22860
rect 21900 21734 22020 22906
rect 22230 22334 22350 22906
rect 22470 21734 22590 22906
rect 22860 21734 22980 22906
rect 25020 22320 25140 22890
rect 25260 22320 25380 22890
rect 26310 22334 26430 22906
rect 26550 21734 26670 22906
rect 26940 21734 27060 22906
rect 27990 22334 28110 22906
rect 28230 21734 28350 22906
rect 28620 21734 28740 22906
rect 29100 22334 29220 22906
rect 29340 22334 29460 22906
rect 29580 22334 29700 22906
rect 30300 21734 30420 22906
rect 30690 21734 30810 22906
rect 30930 22334 31050 22906
rect 31980 22334 32100 22906
rect 32220 22334 32340 22906
rect 32460 22334 32580 22906
rect 33180 22334 33300 22906
rect 33420 22334 33540 22906
rect 33660 22334 33780 22906
rect 34620 22334 34740 22906
rect 34860 22334 34980 22906
rect 35100 22334 35220 22906
rect 35820 22334 35940 22906
rect 36060 22334 36180 22906
rect 36300 22334 36420 22906
rect 36780 21734 36900 22906
rect 37034 21990 37156 22860
rect 37500 21734 37620 22906
rect 37964 21990 38086 22860
rect 38220 21734 38340 22906
rect 39030 22334 39150 22906
rect 39270 21734 39390 22906
rect 39660 21734 39780 22906
rect 40380 22334 40500 22906
rect 40620 22334 40740 22906
rect 40860 22334 40980 22906
rect 41670 22334 41790 22906
rect 41910 21734 42030 22906
rect 42300 21734 42420 22906
rect 43260 21720 43380 22890
rect 43650 21720 43770 22890
rect 44220 21734 44340 22906
rect 44474 21990 44596 22860
rect 44940 21734 45060 22906
rect 45404 21990 45526 22860
rect 45660 21734 45780 22906
rect 45900 21734 46020 22906
rect 46154 21990 46276 22860
rect 46620 21734 46740 22906
rect 47084 21990 47206 22860
rect 47340 21734 47460 22906
rect 47580 22320 47700 22890
rect 47820 22320 47940 22890
rect 48780 21734 48900 22906
rect 49020 21720 49140 22740
rect 49260 21734 49380 22906
rect 49500 21900 49620 22920
rect 49740 21854 49860 22876
rect 5670 17294 5790 17866
rect 5910 17294 6030 18466
rect 6300 17294 6420 18466
rect 8940 17294 9060 18466
rect 9194 17340 9316 18210
rect 9660 17294 9780 18466
rect 10124 17340 10246 18210
rect 10380 17294 10500 18466
rect 11580 17294 11700 18466
rect 11834 17340 11956 18210
rect 12300 17294 12420 18466
rect 12764 17340 12886 18210
rect 13020 17294 13140 18466
rect 13500 17294 13620 18466
rect 13754 17340 13876 18210
rect 14220 17294 14340 18466
rect 14684 17340 14806 18210
rect 14940 17294 15060 18466
rect 15420 17324 15540 18346
rect 15660 17280 15780 18300
rect 15900 17294 16020 18466
rect 16140 17294 16260 18466
rect 17910 17294 18030 17866
rect 18150 17294 18270 18466
rect 18540 17294 18660 18466
rect 19500 17294 19620 17866
rect 19740 17294 19860 17866
rect 19980 17294 20100 17866
rect 20940 17294 21060 17866
rect 21180 17294 21300 17866
rect 21420 17294 21540 17866
rect 22140 17294 22260 17866
rect 22380 17294 22500 17866
rect 22620 17294 22740 17866
rect 23580 17294 23700 17866
rect 23820 17294 23940 17866
rect 24060 17294 24180 17866
rect 24540 17294 24660 18466
rect 24794 17340 24916 18210
rect 25260 17294 25380 18466
rect 25724 17340 25846 18210
rect 25980 17294 26100 18466
rect 26220 17294 26340 18466
rect 26610 17294 26730 18466
rect 26850 17294 26970 17866
rect 27180 17310 27300 17880
rect 27420 17310 27540 17880
rect 28470 17294 28590 17866
rect 28710 17294 28830 18466
rect 29100 17294 29220 18466
rect 30540 17294 30660 17866
rect 30780 17294 30900 17866
rect 31020 17294 31140 17866
rect 31980 17294 32100 17866
rect 32220 17294 32340 17866
rect 32460 17294 32580 17866
rect 33180 17294 33300 18466
rect 33570 17294 33690 18466
rect 33810 17294 33930 17866
rect 35820 17294 35940 17866
rect 36060 17294 36180 17866
rect 36300 17294 36420 17866
rect 36780 17294 36900 18466
rect 37020 17294 37140 18466
rect 37260 17280 37380 18300
rect 37500 17324 37620 18346
rect 37980 17294 38100 17866
rect 38220 17294 38340 17866
rect 38460 17294 38580 17866
rect 38940 17294 39060 17866
rect 39180 17294 39300 17866
rect 39420 17294 39540 17866
rect 40380 17294 40500 17866
rect 40620 17294 40740 17866
rect 40860 17294 40980 17866
rect 41580 17310 41700 17880
rect 41820 17310 41940 17880
rect 42780 17324 42900 18346
rect 43020 17280 43140 18300
rect 43260 17294 43380 18466
rect 43500 17460 43620 18480
rect 43740 17294 43860 18466
rect 44460 17294 44580 18466
rect 44850 17294 44970 18466
rect 45090 17294 45210 17866
rect 46140 17294 46260 17866
rect 46380 17294 46500 17866
rect 46620 17294 46740 17866
rect 47580 17310 47700 18480
rect 47970 17310 48090 18480
rect 49020 17294 49140 18466
rect 49410 17294 49530 18466
rect 49650 17294 49770 17866
rect 6300 16334 6420 16906
rect 6540 16334 6660 16906
rect 6780 16334 6900 16906
rect 7740 15734 7860 16906
rect 7994 15990 8116 16860
rect 8460 15734 8580 16906
rect 8924 15990 9046 16860
rect 9180 15734 9300 16906
rect 9420 15734 9540 16906
rect 9674 15990 9796 16860
rect 10140 15734 10260 16906
rect 10604 15990 10726 16860
rect 10860 15734 10980 16906
rect 11100 15734 11220 16906
rect 11354 15990 11476 16860
rect 11820 15734 11940 16906
rect 12284 15990 12406 16860
rect 12540 15734 12660 16906
rect 13260 15734 13380 16906
rect 13514 15990 13636 16860
rect 13980 15734 14100 16906
rect 14444 15990 14566 16860
rect 14700 15734 14820 16906
rect 14940 15734 15060 16906
rect 15194 15990 15316 16860
rect 15660 15734 15780 16906
rect 16124 15990 16246 16860
rect 16380 15734 16500 16906
rect 16620 15854 16740 16876
rect 16860 15900 16980 16920
rect 17100 15734 17220 16906
rect 17340 15734 17460 16906
rect 17580 16320 17700 16890
rect 17820 16320 17940 16890
rect 18150 16334 18270 16906
rect 18390 15734 18510 16906
rect 18780 15734 18900 16906
rect 19260 16334 19380 16906
rect 19500 16334 19620 16906
rect 19740 16334 19860 16906
rect 20700 15734 20820 16906
rect 21090 15734 21210 16906
rect 21330 16334 21450 16906
rect 22230 16334 22350 16906
rect 22470 15734 22590 16906
rect 22860 15734 22980 16906
rect 23580 16334 23700 16906
rect 23820 16334 23940 16906
rect 24060 16334 24180 16906
rect 24780 16334 24900 16906
rect 25020 16334 25140 16906
rect 25260 16334 25380 16906
rect 25740 15734 25860 16906
rect 25994 15990 26116 16860
rect 26460 15734 26580 16906
rect 26924 15990 27046 16860
rect 27180 15734 27300 16906
rect 27900 16334 28020 16906
rect 28140 16334 28260 16906
rect 28380 16334 28500 16906
rect 29100 16334 29220 16906
rect 29340 16334 29460 16906
rect 29580 16334 29700 16906
rect 30300 15734 30420 16906
rect 30554 15990 30676 16860
rect 31020 15734 31140 16906
rect 31484 15990 31606 16860
rect 31740 15734 31860 16906
rect 32220 16334 32340 16906
rect 32460 16334 32580 16906
rect 32700 16334 32820 16906
rect 33180 16334 33300 16906
rect 33420 16334 33540 16906
rect 33660 16334 33780 16906
rect 34620 16334 34740 16906
rect 34860 16334 34980 16906
rect 35100 16334 35220 16906
rect 36060 15734 36180 16906
rect 36450 15734 36570 16906
rect 36690 16334 36810 16906
rect 37740 16334 37860 16906
rect 37980 16334 38100 16906
rect 38220 16334 38340 16906
rect 38700 15734 38820 16906
rect 38954 15990 39076 16860
rect 39420 15734 39540 16906
rect 39884 15990 40006 16860
rect 40140 15734 40260 16906
rect 41580 15734 41700 16906
rect 41834 15990 41956 16860
rect 42300 15734 42420 16906
rect 42764 15990 42886 16860
rect 43020 15734 43140 16906
rect 44460 15734 44580 16906
rect 44850 15734 44970 16906
rect 45090 16334 45210 16906
rect 46140 16334 46260 16906
rect 46380 16334 46500 16906
rect 46620 16334 46740 16906
rect 47580 16334 47700 16906
rect 47820 16334 47940 16906
rect 48060 16334 48180 16906
rect 49020 15734 49140 16906
rect 49410 15734 49530 16906
rect 49650 16334 49770 16906
rect 6780 11294 6900 11866
rect 7020 11294 7140 11866
rect 7260 11294 7380 11866
rect 8940 11294 9060 12466
rect 9344 11294 9616 12466
rect 9900 11294 10020 12466
rect 10860 11294 10980 11866
rect 11100 11294 11220 11866
rect 11340 11294 11460 11866
rect 12150 11294 12270 11866
rect 12390 11294 12510 12466
rect 12780 11294 12900 12466
rect 15900 11294 16020 11866
rect 16140 11294 16260 11866
rect 16380 11294 16500 11866
rect 16710 11294 16830 11866
rect 16950 11294 17070 12466
rect 17340 11294 17460 12466
rect 17580 11294 17700 12466
rect 17834 11340 17956 12210
rect 18300 11294 18420 12466
rect 18764 11340 18886 12210
rect 19020 11294 19140 12466
rect 19260 11294 19380 12466
rect 19514 11340 19636 12210
rect 19980 11294 20100 12466
rect 20444 11340 20566 12210
rect 20700 11294 20820 12466
rect 21900 11294 22020 12466
rect 22154 11340 22276 12210
rect 22620 11294 22740 12466
rect 23084 11340 23206 12210
rect 23340 11294 23460 12466
rect 25020 11294 25140 12466
rect 25410 11294 25530 12466
rect 25650 11294 25770 11866
rect 26700 11294 26820 11866
rect 26940 11294 27060 11866
rect 27180 11294 27300 11866
rect 29100 11294 29220 12466
rect 29490 11294 29610 12466
rect 29730 11294 29850 11866
rect 30390 11294 30510 11866
rect 30630 11294 30750 12466
rect 31020 11294 31140 12466
rect 31980 11294 32100 11866
rect 32220 11294 32340 11866
rect 32460 11294 32580 11866
rect 32940 11294 33060 12466
rect 33194 11340 33316 12210
rect 33660 11294 33780 12466
rect 34124 11340 34246 12210
rect 34380 11294 34500 12466
rect 34620 11294 34740 12466
rect 35010 11294 35130 12466
rect 35250 11294 35370 11866
rect 36060 11294 36180 11866
rect 36300 11294 36420 11866
rect 36540 11294 36660 11866
rect 37500 11294 37620 11866
rect 37740 11294 37860 11866
rect 37980 11294 38100 11866
rect 38940 11294 39060 11866
rect 39180 11294 39300 11866
rect 39420 11294 39540 11866
rect 40230 11294 40350 11866
rect 40470 11294 40590 12466
rect 40860 11294 40980 12466
rect 41580 11294 41700 11866
rect 41820 11294 41940 11866
rect 42060 11294 42180 11866
rect 42300 11294 42420 11866
rect 43260 11294 43380 11866
rect 43500 11294 43620 11866
rect 43740 11294 43860 11866
rect 44460 11294 44580 12466
rect 44850 11294 44970 12466
rect 45090 11294 45210 11866
rect 46140 11294 46260 11866
rect 46380 11294 46500 11866
rect 46620 11294 46740 11866
rect 47580 11294 47700 12466
rect 47970 11294 48090 12466
rect 48210 11294 48330 11866
rect 49260 11294 49380 11866
rect 49500 11294 49620 11866
rect 49740 11294 49860 11866
rect 5670 10334 5790 10906
rect 5910 9734 6030 10906
rect 6300 9734 6420 10906
rect 6780 10334 6900 10906
rect 7020 10334 7140 10906
rect 7260 10334 7380 10906
rect 7740 9734 7860 10906
rect 7994 9990 8116 10860
rect 8460 9734 8580 10906
rect 8924 9990 9046 10860
rect 9180 9734 9300 10906
rect 9660 10334 9780 10906
rect 9900 10334 10020 10906
rect 10140 10334 10260 10906
rect 10380 10334 10500 10906
rect 11340 10334 11460 10906
rect 11580 10334 11700 10906
rect 11820 10334 11940 10906
rect 13740 9734 13860 10906
rect 13994 9990 14116 10860
rect 14460 9734 14580 10906
rect 14924 9990 15046 10860
rect 15180 9734 15300 10906
rect 16380 10334 16500 10906
rect 16620 10334 16740 10906
rect 16860 10334 16980 10906
rect 17340 9734 17460 10906
rect 17594 9990 17716 10860
rect 18060 9734 18180 10906
rect 18524 9990 18646 10860
rect 18780 9734 18900 10906
rect 19260 9734 19380 10906
rect 19514 9990 19636 10860
rect 19980 9734 20100 10906
rect 20444 9990 20566 10860
rect 20700 9734 20820 10906
rect 21180 10334 21300 10906
rect 21420 10334 21540 10906
rect 21660 10334 21780 10906
rect 21900 9734 22020 10906
rect 22154 9990 22276 10860
rect 22620 9734 22740 10906
rect 23084 9990 23206 10860
rect 23340 9734 23460 10906
rect 23820 10334 23940 10906
rect 24060 10334 24180 10906
rect 24300 10334 24420 10906
rect 25500 9734 25620 10906
rect 25754 9990 25876 10860
rect 26220 9734 26340 10906
rect 26684 9990 26806 10860
rect 26940 9734 27060 10906
rect 27900 10334 28020 10906
rect 28140 10334 28260 10906
rect 28380 10334 28500 10906
rect 29340 10320 29460 10890
rect 29580 10320 29700 10890
rect 30540 10320 30660 10890
rect 30780 10320 30900 10890
rect 31740 9734 31860 10906
rect 32130 9734 32250 10906
rect 32370 10334 32490 10906
rect 33180 9734 33300 10906
rect 33434 9990 33556 10860
rect 33900 9734 34020 10906
rect 34364 9990 34486 10860
rect 34620 9734 34740 10906
rect 35580 10334 35700 10906
rect 35820 10334 35940 10906
rect 36060 10334 36180 10906
rect 36300 10334 36420 10906
rect 36780 10334 36900 10906
rect 37020 10334 37140 10906
rect 37260 10334 37380 10906
rect 37740 10334 37860 10906
rect 37980 10334 38100 10906
rect 38220 10334 38340 10906
rect 38460 10334 38580 10906
rect 38940 9734 39060 10906
rect 39330 9734 39450 10906
rect 39570 10334 39690 10906
rect 40380 10334 40500 10906
rect 40620 10334 40740 10906
rect 40860 10334 40980 10906
rect 41580 10334 41700 10906
rect 41820 10334 41940 10906
rect 42060 10334 42180 10906
rect 42540 9734 42660 10906
rect 42794 9990 42916 10860
rect 43260 9734 43380 10906
rect 43724 9990 43846 10860
rect 43980 9734 44100 10906
rect 45180 9734 45300 10906
rect 45434 9990 45556 10860
rect 45900 9734 46020 10906
rect 46364 9990 46486 10860
rect 46620 9734 46740 10906
rect 47580 10334 47700 10906
rect 47820 10334 47940 10906
rect 48060 10334 48180 10906
rect 49020 10334 49140 10906
rect 49260 10334 49380 10906
rect 49500 10334 49620 10906
rect 5580 5294 5700 6466
rect 5834 5340 5956 6210
rect 6300 5294 6420 6466
rect 6764 5340 6886 6210
rect 7020 5294 7140 6466
rect 7980 5310 8100 5880
rect 8220 5310 8340 5880
rect 8790 5294 8910 5866
rect 9030 5294 9150 6466
rect 9420 5294 9540 6466
rect 9900 5294 10020 5866
rect 10140 5294 10260 5866
rect 10380 5294 10500 5866
rect 10950 5294 11070 5866
rect 11190 5294 11310 6466
rect 11580 5294 11700 6466
rect 12300 5294 12420 5866
rect 12540 5294 12660 5866
rect 12780 5294 12900 5866
rect 13740 5324 13860 6346
rect 13980 5280 14100 6300
rect 14220 5294 14340 6466
rect 14460 5294 14580 6466
rect 15420 5310 15540 6480
rect 15810 5310 15930 6480
rect 18060 5310 18180 6480
rect 18450 5310 18570 6480
rect 20700 5294 20820 5866
rect 20940 5294 21060 5866
rect 21180 5294 21300 5866
rect 23340 5294 23460 5866
rect 23580 5294 23700 5866
rect 23820 5294 23940 5866
rect 25740 5294 25860 6466
rect 25994 5340 26116 6210
rect 26460 5294 26580 6466
rect 26924 5340 27046 6210
rect 27180 5294 27300 6466
rect 27900 5294 28020 5866
rect 28140 5294 28260 5866
rect 28380 5294 28500 5866
rect 29100 5294 29220 5866
rect 29340 5294 29460 5866
rect 29580 5294 29700 5866
rect 30060 5294 30180 6466
rect 30314 5340 30436 6210
rect 30780 5294 30900 6466
rect 31244 5340 31366 6210
rect 31500 5294 31620 6466
rect 31980 5294 32100 6466
rect 32370 5294 32490 6466
rect 32610 5294 32730 5866
rect 33180 5294 33300 5866
rect 33420 5294 33540 5866
rect 33660 5294 33780 5866
rect 34620 5294 34740 5866
rect 34860 5294 34980 5866
rect 35100 5294 35220 5866
rect 36060 5294 36180 5866
rect 36300 5294 36420 5866
rect 36540 5294 36660 5866
rect 37590 5294 37710 5866
rect 37830 5294 37950 6466
rect 38220 5294 38340 6466
rect 38940 5294 39060 5866
rect 39180 5294 39300 5866
rect 39420 5294 39540 5866
rect 40380 5294 40500 5866
rect 40620 5294 40740 5866
rect 40860 5294 40980 5866
rect 43260 5310 43380 6480
rect 43650 5310 43770 6480
rect 44460 5324 44580 6346
rect 44700 5280 44820 6300
rect 44940 5294 45060 6466
rect 45180 5460 45300 6480
rect 45420 5294 45540 6466
rect 46380 5310 46500 5880
rect 46620 5310 46740 5880
rect 47430 5294 47550 5866
rect 47670 5294 47790 6466
rect 48060 5294 48180 6466
<< psubstratepcontact >>
rect 5220 44040 5340 44160
rect 5460 44040 5580 44160
rect 5940 44040 6060 44160
rect 6420 44040 6540 44160
rect 6660 44040 6780 44160
rect 7140 44040 7260 44160
rect 7380 44040 7500 44160
rect 7620 44040 7740 44160
rect 8100 44040 8220 44160
rect 8580 44040 8700 44160
rect 8820 44040 8940 44160
rect 9300 44040 9420 44160
rect 9780 44040 9900 44160
rect 10260 44040 10380 44160
rect 10500 44040 10620 44160
rect 10740 44040 10860 44160
rect 10980 44040 11100 44160
rect 11460 44040 11580 44160
rect 11700 44040 11820 44160
rect 11940 44040 12060 44160
rect 12180 44040 12300 44160
rect 12420 44040 12540 44160
rect 12900 44040 13020 44160
rect 13140 44040 13260 44160
rect 13380 44040 13500 44160
rect 13620 44040 13740 44160
rect 14100 44040 14220 44160
rect 14580 44040 14700 44160
rect 14820 44040 14940 44160
rect 15060 44040 15180 44160
rect 15300 44040 15420 44160
rect 15780 44040 15900 44160
rect 16020 44040 16140 44160
rect 16260 44040 16380 44160
rect 16500 44040 16620 44160
rect 16740 44040 16860 44160
rect 16980 44040 17100 44160
rect 17460 44040 17580 44160
rect 17940 44040 18060 44160
rect 18180 44040 18300 44160
rect 18420 44040 18540 44160
rect 18660 44040 18780 44160
rect 18900 44040 19020 44160
rect 19140 44040 19260 44160
rect 19380 44040 19500 44160
rect 19860 44040 19980 44160
rect 20340 44040 20460 44160
rect 20820 44040 20940 44160
rect 21060 44040 21180 44160
rect 21540 44040 21660 44160
rect 21780 44040 21900 44160
rect 22020 44040 22140 44160
rect 22260 44040 22380 44160
rect 22500 44040 22620 44160
rect 22980 44040 23100 44160
rect 23460 44040 23580 44160
rect 23940 44040 24060 44160
rect 24180 44040 24300 44160
rect 24420 44040 24540 44160
rect 24660 44040 24780 44160
rect 24900 44040 25020 44160
rect 25380 44040 25500 44160
rect 25860 44040 25980 44160
rect 26100 44040 26220 44160
rect 26340 44040 26460 44160
rect 26580 44040 26700 44160
rect 27060 44040 27180 44160
rect 27300 44040 27420 44160
rect 27540 44040 27660 44160
rect 27780 44040 27900 44160
rect 28260 44040 28380 44160
rect 28740 44040 28860 44160
rect 28980 44040 29100 44160
rect 29460 44040 29580 44160
rect 29700 44040 29820 44160
rect 29940 44040 30060 44160
rect 30180 44040 30300 44160
rect 30660 44040 30780 44160
rect 31140 44040 31260 44160
rect 31380 44040 31500 44160
rect 31620 44040 31740 44160
rect 32100 44040 32220 44160
rect 32580 44040 32700 44160
rect 32820 44040 32940 44160
rect 33060 44040 33180 44160
rect 33300 44040 33420 44160
rect 33780 44040 33900 44160
rect 34020 44040 34140 44160
rect 34260 44040 34380 44160
rect 34500 44040 34620 44160
rect 34980 44040 35100 44160
rect 35220 44040 35340 44160
rect 35460 44040 35580 44160
rect 35700 44040 35820 44160
rect 36180 44040 36300 44160
rect 36660 44040 36780 44160
rect 37140 44040 37260 44160
rect 37380 44040 37500 44160
rect 37620 44040 37740 44160
rect 38100 44040 38220 44160
rect 38580 44040 38700 44160
rect 38820 44040 38940 44160
rect 39060 44040 39180 44160
rect 39300 44040 39420 44160
rect 39540 44040 39660 44160
rect 40020 44040 40140 44160
rect 40500 44040 40620 44160
rect 40980 44040 41100 44160
rect 41220 44040 41340 44160
rect 41460 44040 41580 44160
rect 41700 44040 41820 44160
rect 42180 44040 42300 44160
rect 42420 44040 42540 44160
rect 42660 44040 42780 44160
rect 42900 44040 43020 44160
rect 43380 44040 43500 44160
rect 43860 44040 43980 44160
rect 44100 44040 44220 44160
rect 44580 44040 44700 44160
rect 45540 44040 45660 44160
rect 46020 44040 46140 44160
rect 46500 44040 46620 44160
rect 46980 44040 47100 44160
rect 47220 44040 47340 44160
rect 47700 44040 47820 44160
rect 48180 44040 48300 44160
rect 48660 44040 48780 44160
rect 48900 44040 49020 44160
rect 49140 44040 49260 44160
rect 49380 44040 49500 44160
rect 49620 44040 49740 44160
rect 49860 44040 49980 44160
rect 50100 44040 50220 44160
rect 5220 38040 5340 38160
rect 5460 38040 5580 38160
rect 5700 38040 5820 38160
rect 6180 38040 6300 38160
rect 6420 38040 6540 38160
rect 6660 38040 6780 38160
rect 6900 38040 7020 38160
rect 7140 38040 7260 38160
rect 7380 38040 7500 38160
rect 7620 38040 7740 38160
rect 7860 38040 7980 38160
rect 8100 38040 8220 38160
rect 8340 38040 8460 38160
rect 8580 38040 8700 38160
rect 8820 38040 8940 38160
rect 9060 38040 9180 38160
rect 9300 38040 9420 38160
rect 9540 38040 9660 38160
rect 9780 38040 9900 38160
rect 10020 38040 10140 38160
rect 10260 38040 10380 38160
rect 10500 38040 10620 38160
rect 10740 38040 10860 38160
rect 10980 38040 11100 38160
rect 11220 38040 11340 38160
rect 11460 38040 11580 38160
rect 11700 38040 11820 38160
rect 11940 38040 12060 38160
rect 12420 38040 12540 38160
rect 12900 38040 13020 38160
rect 13140 38040 13260 38160
rect 13380 38040 13500 38160
rect 13620 38040 13740 38160
rect 13860 38040 13980 38160
rect 14100 38040 14220 38160
rect 14340 38040 14460 38160
rect 14580 38040 14700 38160
rect 14820 38040 14940 38160
rect 15300 38040 15420 38160
rect 15540 38040 15660 38160
rect 15780 38040 15900 38160
rect 16020 38040 16140 38160
rect 16260 38040 16380 38160
rect 16500 38040 16620 38160
rect 16740 38040 16860 38160
rect 16980 38040 17100 38160
rect 17220 38040 17340 38160
rect 17460 38040 17580 38160
rect 17700 38040 17820 38160
rect 17940 38040 18060 38160
rect 18420 38040 18540 38160
rect 18660 38040 18780 38160
rect 18900 38040 19020 38160
rect 19140 38040 19260 38160
rect 19380 38040 19500 38160
rect 19620 38040 19740 38160
rect 19860 38040 19980 38160
rect 20100 38040 20220 38160
rect 20340 38040 20460 38160
rect 20580 38040 20700 38160
rect 20820 38040 20940 38160
rect 21060 38040 21180 38160
rect 21300 38040 21420 38160
rect 21540 38040 21660 38160
rect 21780 38040 21900 38160
rect 22020 38040 22140 38160
rect 22260 38040 22380 38160
rect 22740 38040 22860 38160
rect 22980 38040 23100 38160
rect 23220 38040 23340 38160
rect 23460 38040 23580 38160
rect 23700 38040 23820 38160
rect 24180 38040 24300 38160
rect 24420 38040 24540 38160
rect 24660 38040 24780 38160
rect 24900 38040 25020 38160
rect 25140 38040 25260 38160
rect 25620 38040 25740 38160
rect 25860 38040 25980 38160
rect 26100 38040 26220 38160
rect 26340 38040 26460 38160
rect 26580 38040 26700 38160
rect 26820 38040 26940 38160
rect 27060 38040 27180 38160
rect 27300 38040 27420 38160
rect 27540 38040 27660 38160
rect 27780 38040 27900 38160
rect 28260 38040 28380 38160
rect 28500 38040 28620 38160
rect 28740 38040 28860 38160
rect 28980 38040 29100 38160
rect 29220 38040 29340 38160
rect 29460 38040 29580 38160
rect 29700 38040 29820 38160
rect 29940 38040 30060 38160
rect 30180 38040 30300 38160
rect 30420 38040 30540 38160
rect 30660 38040 30780 38160
rect 30900 38040 31020 38160
rect 31140 38040 31260 38160
rect 31380 38040 31500 38160
rect 31620 38040 31740 38160
rect 31860 38040 31980 38160
rect 32100 38040 32220 38160
rect 32340 38040 32460 38160
rect 32580 38040 32700 38160
rect 32820 38040 32940 38160
rect 33060 38040 33180 38160
rect 33300 38040 33420 38160
rect 33780 38040 33900 38160
rect 34020 38040 34140 38160
rect 34260 38040 34380 38160
rect 34500 38040 34620 38160
rect 34740 38040 34860 38160
rect 34980 38040 35100 38160
rect 35220 38040 35340 38160
rect 35460 38040 35580 38160
rect 35700 38040 35820 38160
rect 35940 38040 36060 38160
rect 36180 38040 36300 38160
rect 36420 38040 36540 38160
rect 36660 38040 36780 38160
rect 36900 38040 37020 38160
rect 37140 38040 37260 38160
rect 37380 38040 37500 38160
rect 37620 38040 37740 38160
rect 37860 38040 37980 38160
rect 38100 38040 38220 38160
rect 38340 38040 38460 38160
rect 38580 38040 38700 38160
rect 38820 38040 38940 38160
rect 39300 38040 39420 38160
rect 39540 38040 39660 38160
rect 39780 38040 39900 38160
rect 40020 38040 40140 38160
rect 40260 38040 40380 38160
rect 40500 38040 40620 38160
rect 40740 38040 40860 38160
rect 40980 38040 41100 38160
rect 41220 38040 41340 38160
rect 41460 38040 41580 38160
rect 41700 38040 41820 38160
rect 41940 38040 42060 38160
rect 42180 38040 42300 38160
rect 42420 38040 42540 38160
rect 42660 38040 42780 38160
rect 42900 38040 43020 38160
rect 43140 38040 43260 38160
rect 43380 38040 43500 38160
rect 43860 38040 43980 38160
rect 44100 38040 44220 38160
rect 44340 38040 44460 38160
rect 44580 38040 44700 38160
rect 44820 38040 44940 38160
rect 45060 38040 45180 38160
rect 45300 38040 45420 38160
rect 45540 38040 45660 38160
rect 45780 38040 45900 38160
rect 46020 38040 46140 38160
rect 46260 38040 46380 38160
rect 46500 38040 46620 38160
rect 46740 38040 46860 38160
rect 46980 38040 47100 38160
rect 47220 38040 47340 38160
rect 47460 38040 47580 38160
rect 47940 38040 48060 38160
rect 48420 38040 48540 38160
rect 48660 38040 48780 38160
rect 48900 38040 49020 38160
rect 49140 38040 49260 38160
rect 49380 38040 49500 38160
rect 49860 38040 49980 38160
rect 50100 38040 50220 38160
rect 5220 32040 5340 32160
rect 5460 32040 5580 32160
rect 5700 32040 5820 32160
rect 5940 32040 6060 32160
rect 6180 32040 6300 32160
rect 6420 32040 6540 32160
rect 6900 32040 7020 32160
rect 7140 32040 7260 32160
rect 7380 32040 7500 32160
rect 7620 32040 7740 32160
rect 7860 32040 7980 32160
rect 8100 32040 8220 32160
rect 8340 32040 8460 32160
rect 8580 32040 8700 32160
rect 8820 32040 8940 32160
rect 9060 32040 9180 32160
rect 9300 32040 9420 32160
rect 9540 32040 9660 32160
rect 9780 32040 9900 32160
rect 10260 32040 10380 32160
rect 10500 32040 10620 32160
rect 10740 32040 10860 32160
rect 10980 32040 11100 32160
rect 11460 32040 11580 32160
rect 11940 32040 12060 32160
rect 12420 32040 12540 32160
rect 12660 32040 12780 32160
rect 12900 32040 13020 32160
rect 13140 32040 13260 32160
rect 13380 32040 13500 32160
rect 13620 32040 13740 32160
rect 13860 32040 13980 32160
rect 14100 32040 14220 32160
rect 14340 32040 14460 32160
rect 14580 32040 14700 32160
rect 14820 32040 14940 32160
rect 15060 32040 15180 32160
rect 15540 32040 15660 32160
rect 15780 32040 15900 32160
rect 16020 32040 16140 32160
rect 16260 32040 16380 32160
rect 16500 32040 16620 32160
rect 16740 32040 16860 32160
rect 16980 32040 17100 32160
rect 17460 32040 17580 32160
rect 17700 32040 17820 32160
rect 17940 32040 18060 32160
rect 18180 32040 18300 32160
rect 18420 32040 18540 32160
rect 18660 32040 18780 32160
rect 18900 32040 19020 32160
rect 19140 32040 19260 32160
rect 19380 32040 19500 32160
rect 19620 32040 19740 32160
rect 19860 32040 19980 32160
rect 20100 32040 20220 32160
rect 20340 32040 20460 32160
rect 20580 32040 20700 32160
rect 20820 32040 20940 32160
rect 21060 32040 21180 32160
rect 21540 32040 21660 32160
rect 21780 32040 21900 32160
rect 22020 32040 22140 32160
rect 22260 32040 22380 32160
rect 22500 32040 22620 32160
rect 22740 32040 22860 32160
rect 22980 32040 23100 32160
rect 23220 32040 23340 32160
rect 23460 32040 23580 32160
rect 23700 32040 23820 32160
rect 24180 32040 24300 32160
rect 24420 32040 24540 32160
rect 24660 32040 24780 32160
rect 25140 32040 25260 32160
rect 25620 32040 25740 32160
rect 25860 32040 25980 32160
rect 26340 32040 26460 32160
rect 26820 32040 26940 32160
rect 27060 32040 27180 32160
rect 27300 32040 27420 32160
rect 27540 32040 27660 32160
rect 27780 32040 27900 32160
rect 28020 32040 28140 32160
rect 28260 32040 28380 32160
rect 28500 32040 28620 32160
rect 28740 32040 28860 32160
rect 28980 32040 29100 32160
rect 29220 32040 29340 32160
rect 29460 32040 29580 32160
rect 29700 32040 29820 32160
rect 29940 32040 30060 32160
rect 30180 32040 30300 32160
rect 30420 32040 30540 32160
rect 30660 32040 30780 32160
rect 30900 32040 31020 32160
rect 31140 32040 31260 32160
rect 31380 32040 31500 32160
rect 31620 32040 31740 32160
rect 31860 32040 31980 32160
rect 32340 32040 32460 32160
rect 32580 32040 32700 32160
rect 32820 32040 32940 32160
rect 33060 32040 33180 32160
rect 33540 32040 33660 32160
rect 33780 32040 33900 32160
rect 34020 32040 34140 32160
rect 34260 32040 34380 32160
rect 34500 32040 34620 32160
rect 34980 32040 35100 32160
rect 35220 32040 35340 32160
rect 35460 32040 35580 32160
rect 35700 32040 35820 32160
rect 35940 32040 36060 32160
rect 36420 32040 36540 32160
rect 36660 32040 36780 32160
rect 36900 32040 37020 32160
rect 37140 32040 37260 32160
rect 37380 32040 37500 32160
rect 37620 32040 37740 32160
rect 38100 32040 38220 32160
rect 38340 32040 38460 32160
rect 38580 32040 38700 32160
rect 38820 32040 38940 32160
rect 39300 32040 39420 32160
rect 39540 32040 39660 32160
rect 39780 32040 39900 32160
rect 40020 32040 40140 32160
rect 40260 32040 40380 32160
rect 40500 32040 40620 32160
rect 40980 32040 41100 32160
rect 41220 32040 41340 32160
rect 41460 32040 41580 32160
rect 41700 32040 41820 32160
rect 41940 32040 42060 32160
rect 42180 32040 42300 32160
rect 42420 32040 42540 32160
rect 42660 32040 42780 32160
rect 42900 32040 43020 32160
rect 43380 32040 43500 32160
rect 43860 32040 43980 32160
rect 44100 32040 44220 32160
rect 44340 32040 44460 32160
rect 44580 32040 44700 32160
rect 44820 32040 44940 32160
rect 45060 32040 45180 32160
rect 45300 32040 45420 32160
rect 45540 32040 45660 32160
rect 45780 32040 45900 32160
rect 46020 32040 46140 32160
rect 46260 32040 46380 32160
rect 46500 32040 46620 32160
rect 46740 32040 46860 32160
rect 46980 32040 47100 32160
rect 47220 32040 47340 32160
rect 47460 32040 47580 32160
rect 47700 32040 47820 32160
rect 47940 32040 48060 32160
rect 48180 32040 48300 32160
rect 48420 32040 48540 32160
rect 48660 32040 48780 32160
rect 48900 32040 49020 32160
rect 49140 32040 49260 32160
rect 49380 32040 49500 32160
rect 49620 32040 49740 32160
rect 49860 32040 49980 32160
rect 50100 32040 50220 32160
rect 5220 26040 5340 26160
rect 5460 26040 5580 26160
rect 5700 26040 5820 26160
rect 5940 26040 6060 26160
rect 6180 26040 6300 26160
rect 6420 26040 6540 26160
rect 6660 26040 6780 26160
rect 6900 26040 7020 26160
rect 7380 26040 7500 26160
rect 7860 26040 7980 26160
rect 8100 26040 8220 26160
rect 8340 26040 8460 26160
rect 8580 26040 8700 26160
rect 9060 26040 9180 26160
rect 9300 26040 9420 26160
rect 9540 26040 9660 26160
rect 9780 26040 9900 26160
rect 10020 26040 10140 26160
rect 10260 26040 10380 26160
rect 10500 26040 10620 26160
rect 10740 26040 10860 26160
rect 10980 26040 11100 26160
rect 11220 26040 11340 26160
rect 11460 26040 11580 26160
rect 11700 26040 11820 26160
rect 11940 26040 12060 26160
rect 12420 26040 12540 26160
rect 12660 26040 12780 26160
rect 12900 26040 13020 26160
rect 13140 26040 13260 26160
rect 13380 26040 13500 26160
rect 13620 26040 13740 26160
rect 14100 26040 14220 26160
rect 14340 26040 14460 26160
rect 14580 26040 14700 26160
rect 14820 26040 14940 26160
rect 15060 26040 15180 26160
rect 15300 26040 15420 26160
rect 15780 26040 15900 26160
rect 16020 26040 16140 26160
rect 16260 26040 16380 26160
rect 16500 26040 16620 26160
rect 16740 26040 16860 26160
rect 16980 26040 17100 26160
rect 17220 26040 17340 26160
rect 17460 26040 17580 26160
rect 17700 26040 17820 26160
rect 17940 26040 18060 26160
rect 18180 26040 18300 26160
rect 18420 26040 18540 26160
rect 18660 26040 18780 26160
rect 18900 26040 19020 26160
rect 19140 26040 19260 26160
rect 19380 26040 19500 26160
rect 19620 26040 19740 26160
rect 19860 26040 19980 26160
rect 20100 26040 20220 26160
rect 20340 26040 20460 26160
rect 20580 26040 20700 26160
rect 20820 26040 20940 26160
rect 21300 26040 21420 26160
rect 21540 26040 21660 26160
rect 21780 26040 21900 26160
rect 22020 26040 22140 26160
rect 22260 26040 22380 26160
rect 22500 26040 22620 26160
rect 22740 26040 22860 26160
rect 22980 26040 23100 26160
rect 23220 26040 23340 26160
rect 23460 26040 23580 26160
rect 23700 26040 23820 26160
rect 23940 26040 24060 26160
rect 24180 26040 24300 26160
rect 24420 26040 24540 26160
rect 24660 26040 24780 26160
rect 24900 26040 25020 26160
rect 25140 26040 25260 26160
rect 25380 26040 25500 26160
rect 25620 26040 25740 26160
rect 25860 26040 25980 26160
rect 26100 26040 26220 26160
rect 26340 26040 26460 26160
rect 26580 26040 26700 26160
rect 26820 26040 26940 26160
rect 27060 26040 27180 26160
rect 27300 26040 27420 26160
rect 27540 26040 27660 26160
rect 27780 26040 27900 26160
rect 28020 26040 28140 26160
rect 28260 26040 28380 26160
rect 28740 26040 28860 26160
rect 28980 26040 29100 26160
rect 29220 26040 29340 26160
rect 29460 26040 29580 26160
rect 29700 26040 29820 26160
rect 29940 26040 30060 26160
rect 30180 26040 30300 26160
rect 30420 26040 30540 26160
rect 30660 26040 30780 26160
rect 30900 26040 31020 26160
rect 31140 26040 31260 26160
rect 31380 26040 31500 26160
rect 31620 26040 31740 26160
rect 31860 26040 31980 26160
rect 32100 26040 32220 26160
rect 32580 26040 32700 26160
rect 32820 26040 32940 26160
rect 33060 26040 33180 26160
rect 33300 26040 33420 26160
rect 33540 26040 33660 26160
rect 33780 26040 33900 26160
rect 34020 26040 34140 26160
rect 34260 26040 34380 26160
rect 34500 26040 34620 26160
rect 34740 26040 34860 26160
rect 34980 26040 35100 26160
rect 35220 26040 35340 26160
rect 35460 26040 35580 26160
rect 35700 26040 35820 26160
rect 35940 26040 36060 26160
rect 36420 26040 36540 26160
rect 36660 26040 36780 26160
rect 36900 26040 37020 26160
rect 37140 26040 37260 26160
rect 37380 26040 37500 26160
rect 37620 26040 37740 26160
rect 37860 26040 37980 26160
rect 38100 26040 38220 26160
rect 38340 26040 38460 26160
rect 38580 26040 38700 26160
rect 38820 26040 38940 26160
rect 39060 26040 39180 26160
rect 39300 26040 39420 26160
rect 39540 26040 39660 26160
rect 39780 26040 39900 26160
rect 40020 26040 40140 26160
rect 40260 26040 40380 26160
rect 40500 26040 40620 26160
rect 40740 26040 40860 26160
rect 40980 26040 41100 26160
rect 41220 26040 41340 26160
rect 41460 26040 41580 26160
rect 41700 26040 41820 26160
rect 41940 26040 42060 26160
rect 42180 26040 42300 26160
rect 42420 26040 42540 26160
rect 42660 26040 42780 26160
rect 42900 26040 43020 26160
rect 43140 26040 43260 26160
rect 43380 26040 43500 26160
rect 43620 26040 43740 26160
rect 43860 26040 43980 26160
rect 44100 26040 44220 26160
rect 44340 26040 44460 26160
rect 44820 26040 44940 26160
rect 45060 26040 45180 26160
rect 45300 26040 45420 26160
rect 45540 26040 45660 26160
rect 45780 26040 45900 26160
rect 46020 26040 46140 26160
rect 46260 26040 46380 26160
rect 46500 26040 46620 26160
rect 46740 26040 46860 26160
rect 46980 26040 47100 26160
rect 47220 26040 47340 26160
rect 47460 26040 47580 26160
rect 47700 26040 47820 26160
rect 47940 26040 48060 26160
rect 48180 26040 48300 26160
rect 48420 26040 48540 26160
rect 48660 26040 48780 26160
rect 48900 26040 49020 26160
rect 49140 26040 49260 26160
rect 49380 26040 49500 26160
rect 49620 26040 49740 26160
rect 49860 26040 49980 26160
rect 50100 26040 50220 26160
rect 5220 20040 5340 20160
rect 5460 20040 5580 20160
rect 5700 20040 5820 20160
rect 5940 20040 6060 20160
rect 6180 20040 6300 20160
rect 6420 20040 6540 20160
rect 6660 20040 6780 20160
rect 6900 20040 7020 20160
rect 7140 20040 7260 20160
rect 7380 20040 7500 20160
rect 7620 20040 7740 20160
rect 7860 20040 7980 20160
rect 8100 20040 8220 20160
rect 8340 20040 8460 20160
rect 8580 20040 8700 20160
rect 8820 20040 8940 20160
rect 9060 20040 9180 20160
rect 9300 20040 9420 20160
rect 9540 20040 9660 20160
rect 10020 20040 10140 20160
rect 10260 20040 10380 20160
rect 10500 20040 10620 20160
rect 10740 20040 10860 20160
rect 10980 20040 11100 20160
rect 11220 20040 11340 20160
rect 11460 20040 11580 20160
rect 11940 20040 12060 20160
rect 12180 20040 12300 20160
rect 12420 20040 12540 20160
rect 12660 20040 12780 20160
rect 12900 20040 13020 20160
rect 13140 20040 13260 20160
rect 13380 20040 13500 20160
rect 13620 20040 13740 20160
rect 13860 20040 13980 20160
rect 14100 20040 14220 20160
rect 14340 20040 14460 20160
rect 14580 20040 14700 20160
rect 14820 20040 14940 20160
rect 15060 20040 15180 20160
rect 15300 20040 15420 20160
rect 15540 20040 15660 20160
rect 15780 20040 15900 20160
rect 16020 20040 16140 20160
rect 16260 20040 16380 20160
rect 16500 20040 16620 20160
rect 16740 20040 16860 20160
rect 16980 20040 17100 20160
rect 17220 20040 17340 20160
rect 17460 20040 17580 20160
rect 17700 20040 17820 20160
rect 17940 20040 18060 20160
rect 18180 20040 18300 20160
rect 18420 20040 18540 20160
rect 18660 20040 18780 20160
rect 18900 20040 19020 20160
rect 19140 20040 19260 20160
rect 19380 20040 19500 20160
rect 19860 20040 19980 20160
rect 20100 20040 20220 20160
rect 20340 20040 20460 20160
rect 20580 20040 20700 20160
rect 20820 20040 20940 20160
rect 21060 20040 21180 20160
rect 21300 20040 21420 20160
rect 21540 20040 21660 20160
rect 21780 20040 21900 20160
rect 22020 20040 22140 20160
rect 22500 20040 22620 20160
rect 22740 20040 22860 20160
rect 22980 20040 23100 20160
rect 23220 20040 23340 20160
rect 23460 20040 23580 20160
rect 23700 20040 23820 20160
rect 23940 20040 24060 20160
rect 24180 20040 24300 20160
rect 24420 20040 24540 20160
rect 24660 20040 24780 20160
rect 24900 20040 25020 20160
rect 25380 20040 25500 20160
rect 25620 20040 25740 20160
rect 25860 20040 25980 20160
rect 26100 20040 26220 20160
rect 26580 20040 26700 20160
rect 27060 20040 27180 20160
rect 27300 20040 27420 20160
rect 27540 20040 27660 20160
rect 27780 20040 27900 20160
rect 28020 20040 28140 20160
rect 28260 20040 28380 20160
rect 28740 20040 28860 20160
rect 28980 20040 29100 20160
rect 29220 20040 29340 20160
rect 29460 20040 29580 20160
rect 29700 20040 29820 20160
rect 29940 20040 30060 20160
rect 30180 20040 30300 20160
rect 30420 20040 30540 20160
rect 30660 20040 30780 20160
rect 30900 20040 31020 20160
rect 31140 20040 31260 20160
rect 31380 20040 31500 20160
rect 31620 20040 31740 20160
rect 31860 20040 31980 20160
rect 32340 20040 32460 20160
rect 32580 20040 32700 20160
rect 32820 20040 32940 20160
rect 33060 20040 33180 20160
rect 33540 20040 33660 20160
rect 33780 20040 33900 20160
rect 34020 20040 34140 20160
rect 34260 20040 34380 20160
rect 34500 20040 34620 20160
rect 34740 20040 34860 20160
rect 34980 20040 35100 20160
rect 35220 20040 35340 20160
rect 35460 20040 35580 20160
rect 35700 20040 35820 20160
rect 36180 20040 36300 20160
rect 36420 20040 36540 20160
rect 36660 20040 36780 20160
rect 37140 20040 37260 20160
rect 37620 20040 37740 20160
rect 37860 20040 37980 20160
rect 38100 20040 38220 20160
rect 38340 20040 38460 20160
rect 38580 20040 38700 20160
rect 38820 20040 38940 20160
rect 39300 20040 39420 20160
rect 39540 20040 39660 20160
rect 39780 20040 39900 20160
rect 40020 20040 40140 20160
rect 40260 20040 40380 20160
rect 40740 20040 40860 20160
rect 40980 20040 41100 20160
rect 41220 20040 41340 20160
rect 41460 20040 41580 20160
rect 41940 20040 42060 20160
rect 42180 20040 42300 20160
rect 42420 20040 42540 20160
rect 42660 20040 42780 20160
rect 42900 20040 43020 20160
rect 43140 20040 43260 20160
rect 43620 20040 43740 20160
rect 43860 20040 43980 20160
rect 44100 20040 44220 20160
rect 44340 20040 44460 20160
rect 44580 20040 44700 20160
rect 44820 20040 44940 20160
rect 45060 20040 45180 20160
rect 45300 20040 45420 20160
rect 45540 20040 45660 20160
rect 45780 20040 45900 20160
rect 46020 20040 46140 20160
rect 46500 20040 46620 20160
rect 46740 20040 46860 20160
rect 46980 20040 47100 20160
rect 47220 20040 47340 20160
rect 47460 20040 47580 20160
rect 47940 20040 48060 20160
rect 48180 20040 48300 20160
rect 48420 20040 48540 20160
rect 48660 20040 48780 20160
rect 48900 20040 49020 20160
rect 49380 20040 49500 20160
rect 49860 20040 49980 20160
rect 50100 20040 50220 20160
rect 5220 14040 5340 14160
rect 5460 14040 5580 14160
rect 5700 14040 5820 14160
rect 5940 14040 6060 14160
rect 6180 14040 6300 14160
rect 6420 14040 6540 14160
rect 6660 14040 6780 14160
rect 6900 14040 7020 14160
rect 7140 14040 7260 14160
rect 7380 14040 7500 14160
rect 7620 14040 7740 14160
rect 7860 14040 7980 14160
rect 8100 14040 8220 14160
rect 8340 14040 8460 14160
rect 8580 14040 8700 14160
rect 8820 14040 8940 14160
rect 9060 14040 9180 14160
rect 9300 14040 9420 14160
rect 9780 14040 9900 14160
rect 10020 14040 10140 14160
rect 10260 14040 10380 14160
rect 10500 14040 10620 14160
rect 10740 14040 10860 14160
rect 10980 14040 11100 14160
rect 11220 14040 11340 14160
rect 11460 14040 11580 14160
rect 11700 14040 11820 14160
rect 11940 14040 12060 14160
rect 12420 14040 12540 14160
rect 12660 14040 12780 14160
rect 12900 14040 13020 14160
rect 13140 14040 13260 14160
rect 13380 14040 13500 14160
rect 13620 14040 13740 14160
rect 13860 14040 13980 14160
rect 14100 14040 14220 14160
rect 14340 14040 14460 14160
rect 14580 14040 14700 14160
rect 14820 14040 14940 14160
rect 15060 14040 15180 14160
rect 15300 14040 15420 14160
rect 15540 14040 15660 14160
rect 15780 14040 15900 14160
rect 16260 14040 16380 14160
rect 16500 14040 16620 14160
rect 16980 14040 17100 14160
rect 17460 14040 17580 14160
rect 17940 14040 18060 14160
rect 18420 14040 18540 14160
rect 18900 14040 19020 14160
rect 19140 14040 19260 14160
rect 19380 14040 19500 14160
rect 19620 14040 19740 14160
rect 19860 14040 19980 14160
rect 20100 14040 20220 14160
rect 20340 14040 20460 14160
rect 20580 14040 20700 14160
rect 20820 14040 20940 14160
rect 21060 14040 21180 14160
rect 21300 14040 21420 14160
rect 21540 14040 21660 14160
rect 21780 14040 21900 14160
rect 22020 14040 22140 14160
rect 22260 14040 22380 14160
rect 22500 14040 22620 14160
rect 22740 14040 22860 14160
rect 22980 14040 23100 14160
rect 23220 14040 23340 14160
rect 23460 14040 23580 14160
rect 23700 14040 23820 14160
rect 23940 14040 24060 14160
rect 24180 14040 24300 14160
rect 24420 14040 24540 14160
rect 24660 14040 24780 14160
rect 24900 14040 25020 14160
rect 25380 14040 25500 14160
rect 25620 14040 25740 14160
rect 25860 14040 25980 14160
rect 26100 14040 26220 14160
rect 26340 14040 26460 14160
rect 26580 14040 26700 14160
rect 26820 14040 26940 14160
rect 27060 14040 27180 14160
rect 27300 14040 27420 14160
rect 27540 14040 27660 14160
rect 27780 14040 27900 14160
rect 28020 14040 28140 14160
rect 28260 14040 28380 14160
rect 28500 14040 28620 14160
rect 28740 14040 28860 14160
rect 28980 14040 29100 14160
rect 29460 14040 29580 14160
rect 29700 14040 29820 14160
rect 29940 14040 30060 14160
rect 30180 14040 30300 14160
rect 30420 14040 30540 14160
rect 30660 14040 30780 14160
rect 30900 14040 31020 14160
rect 31140 14040 31260 14160
rect 31380 14040 31500 14160
rect 31620 14040 31740 14160
rect 31860 14040 31980 14160
rect 32100 14040 32220 14160
rect 32340 14040 32460 14160
rect 32580 14040 32700 14160
rect 32820 14040 32940 14160
rect 33060 14040 33180 14160
rect 33300 14040 33420 14160
rect 33540 14040 33660 14160
rect 33780 14040 33900 14160
rect 34020 14040 34140 14160
rect 34260 14040 34380 14160
rect 34500 14040 34620 14160
rect 34980 14040 35100 14160
rect 35220 14040 35340 14160
rect 35460 14040 35580 14160
rect 35700 14040 35820 14160
rect 35940 14040 36060 14160
rect 36420 14040 36540 14160
rect 36660 14040 36780 14160
rect 36900 14040 37020 14160
rect 37140 14040 37260 14160
rect 37380 14040 37500 14160
rect 37620 14040 37740 14160
rect 37860 14040 37980 14160
rect 38100 14040 38220 14160
rect 38340 14040 38460 14160
rect 38580 14040 38700 14160
rect 38820 14040 38940 14160
rect 39300 14040 39420 14160
rect 39540 14040 39660 14160
rect 39780 14040 39900 14160
rect 40020 14040 40140 14160
rect 40260 14040 40380 14160
rect 40500 14040 40620 14160
rect 40740 14040 40860 14160
rect 40980 14040 41100 14160
rect 41220 14040 41340 14160
rect 41460 14040 41580 14160
rect 41940 14040 42060 14160
rect 42420 14040 42540 14160
rect 42660 14040 42780 14160
rect 42900 14040 43020 14160
rect 43140 14040 43260 14160
rect 43380 14040 43500 14160
rect 43620 14040 43740 14160
rect 43860 14040 43980 14160
rect 44100 14040 44220 14160
rect 44340 14040 44460 14160
rect 44820 14040 44940 14160
rect 45300 14040 45420 14160
rect 45540 14040 45660 14160
rect 45780 14040 45900 14160
rect 46020 14040 46140 14160
rect 46500 14040 46620 14160
rect 46740 14040 46860 14160
rect 46980 14040 47100 14160
rect 47220 14040 47340 14160
rect 47460 14040 47580 14160
rect 47700 14040 47820 14160
rect 47940 14040 48060 14160
rect 48180 14040 48300 14160
rect 48420 14040 48540 14160
rect 48660 14040 48780 14160
rect 48900 14040 49020 14160
rect 49140 14040 49260 14160
rect 49380 14040 49500 14160
rect 49860 14040 49980 14160
rect 50100 14040 50220 14160
rect 5220 8040 5340 8160
rect 5460 8040 5580 8160
rect 5700 8040 5820 8160
rect 5940 8040 6060 8160
rect 6180 8040 6300 8160
rect 6420 8040 6540 8160
rect 6660 8040 6780 8160
rect 7140 8040 7260 8160
rect 7380 8040 7500 8160
rect 7620 8040 7740 8160
rect 7860 8040 7980 8160
rect 8100 8040 8220 8160
rect 8340 8040 8460 8160
rect 8580 8040 8700 8160
rect 9060 8040 9180 8160
rect 9300 8040 9420 8160
rect 9540 8040 9660 8160
rect 9780 8040 9900 8160
rect 10020 8040 10140 8160
rect 10260 8040 10380 8160
rect 10500 8040 10620 8160
rect 10740 8040 10860 8160
rect 10980 8040 11100 8160
rect 11220 8040 11340 8160
rect 11460 8040 11580 8160
rect 11700 8040 11820 8160
rect 11940 8040 12060 8160
rect 12180 8040 12300 8160
rect 12420 8040 12540 8160
rect 12660 8040 12780 8160
rect 12900 8040 13020 8160
rect 13140 8040 13260 8160
rect 13380 8040 13500 8160
rect 13620 8040 13740 8160
rect 14100 8040 14220 8160
rect 14580 8040 14700 8160
rect 14820 8040 14940 8160
rect 15060 8040 15180 8160
rect 15300 8040 15420 8160
rect 15540 8040 15660 8160
rect 15780 8040 15900 8160
rect 16020 8040 16140 8160
rect 16260 8040 16380 8160
rect 16500 8040 16620 8160
rect 16740 8040 16860 8160
rect 16980 8040 17100 8160
rect 17220 8040 17340 8160
rect 17460 8040 17580 8160
rect 17700 8040 17820 8160
rect 17940 8040 18060 8160
rect 18180 8040 18300 8160
rect 18420 8040 18540 8160
rect 18660 8040 18780 8160
rect 18900 8040 19020 8160
rect 19140 8040 19260 8160
rect 19380 8040 19500 8160
rect 19620 8040 19740 8160
rect 19860 8040 19980 8160
rect 20100 8040 20220 8160
rect 20340 8040 20460 8160
rect 20580 8040 20700 8160
rect 20820 8040 20940 8160
rect 21060 8040 21180 8160
rect 21300 8040 21420 8160
rect 21540 8040 21660 8160
rect 21780 8040 21900 8160
rect 22020 8040 22140 8160
rect 22260 8040 22380 8160
rect 22500 8040 22620 8160
rect 22740 8040 22860 8160
rect 22980 8040 23100 8160
rect 23220 8040 23340 8160
rect 23460 8040 23580 8160
rect 23700 8040 23820 8160
rect 23940 8040 24060 8160
rect 24180 8040 24300 8160
rect 24420 8040 24540 8160
rect 24660 8040 24780 8160
rect 24900 8040 25020 8160
rect 25140 8040 25260 8160
rect 25380 8040 25500 8160
rect 25620 8040 25740 8160
rect 25860 8040 25980 8160
rect 26100 8040 26220 8160
rect 26340 8040 26460 8160
rect 26580 8040 26700 8160
rect 26820 8040 26940 8160
rect 27060 8040 27180 8160
rect 27300 8040 27420 8160
rect 27540 8040 27660 8160
rect 27780 8040 27900 8160
rect 28260 8040 28380 8160
rect 28500 8040 28620 8160
rect 28740 8040 28860 8160
rect 28980 8040 29100 8160
rect 29220 8040 29340 8160
rect 29460 8040 29580 8160
rect 29700 8040 29820 8160
rect 29940 8040 30060 8160
rect 30180 8040 30300 8160
rect 30420 8040 30540 8160
rect 30900 8040 31020 8160
rect 31140 8040 31260 8160
rect 31380 8040 31500 8160
rect 31620 8040 31740 8160
rect 31860 8040 31980 8160
rect 32100 8040 32220 8160
rect 32340 8040 32460 8160
rect 32580 8040 32700 8160
rect 32820 8040 32940 8160
rect 33060 8040 33180 8160
rect 33300 8040 33420 8160
rect 33540 8040 33660 8160
rect 33780 8040 33900 8160
rect 34020 8040 34140 8160
rect 34260 8040 34380 8160
rect 34500 8040 34620 8160
rect 34740 8040 34860 8160
rect 34980 8040 35100 8160
rect 35220 8040 35340 8160
rect 35460 8040 35580 8160
rect 35700 8040 35820 8160
rect 35940 8040 36060 8160
rect 36420 8040 36540 8160
rect 36660 8040 36780 8160
rect 36900 8040 37020 8160
rect 37140 8040 37260 8160
rect 37380 8040 37500 8160
rect 37620 8040 37740 8160
rect 37860 8040 37980 8160
rect 38100 8040 38220 8160
rect 38340 8040 38460 8160
rect 38580 8040 38700 8160
rect 38820 8040 38940 8160
rect 39300 8040 39420 8160
rect 39540 8040 39660 8160
rect 39780 8040 39900 8160
rect 40020 8040 40140 8160
rect 40260 8040 40380 8160
rect 40740 8040 40860 8160
rect 40980 8040 41100 8160
rect 41220 8040 41340 8160
rect 41460 8040 41580 8160
rect 41700 8040 41820 8160
rect 41940 8040 42060 8160
rect 42180 8040 42300 8160
rect 42420 8040 42540 8160
rect 42660 8040 42780 8160
rect 42900 8040 43020 8160
rect 43140 8040 43260 8160
rect 43380 8040 43500 8160
rect 43620 8040 43740 8160
rect 43860 8040 43980 8160
rect 44100 8040 44220 8160
rect 44340 8040 44460 8160
rect 44580 8040 44700 8160
rect 44820 8040 44940 8160
rect 45060 8040 45180 8160
rect 45300 8040 45420 8160
rect 45540 8040 45660 8160
rect 45780 8040 45900 8160
rect 46020 8040 46140 8160
rect 46260 8040 46380 8160
rect 46500 8040 46620 8160
rect 46740 8040 46860 8160
rect 46980 8040 47100 8160
rect 47220 8040 47340 8160
rect 47460 8040 47580 8160
rect 47700 8040 47820 8160
rect 48180 8040 48300 8160
rect 48420 8040 48540 8160
rect 48660 8040 48780 8160
rect 48900 8040 49020 8160
rect 49140 8040 49260 8160
rect 49380 8040 49500 8160
rect 49620 8040 49740 8160
rect 49860 8040 49980 8160
rect 50100 8040 50220 8160
<< nsubstratencontact >>
rect 5220 41040 5340 41160
rect 5460 41040 5580 41160
rect 5700 41040 5820 41160
rect 5940 41040 6060 41160
rect 6180 41040 6300 41160
rect 6420 41040 6540 41160
rect 6660 41040 6780 41160
rect 6900 41040 7020 41160
rect 7140 41040 7260 41160
rect 7380 41040 7500 41160
rect 7620 41040 7740 41160
rect 7860 41040 7980 41160
rect 8100 41040 8220 41160
rect 8340 41040 8460 41160
rect 8580 41040 8700 41160
rect 8820 41040 8940 41160
rect 9060 41040 9180 41160
rect 9300 41040 9420 41160
rect 9540 41040 9660 41160
rect 9780 41040 9900 41160
rect 10020 41040 10140 41160
rect 10260 41040 10380 41160
rect 10500 41040 10620 41160
rect 10740 41040 10860 41160
rect 10980 41040 11100 41160
rect 11460 41040 11580 41160
rect 11700 41040 11820 41160
rect 11940 41040 12060 41160
rect 12180 41040 12300 41160
rect 12420 41040 12540 41160
rect 12900 41040 13020 41160
rect 13140 41040 13260 41160
rect 13380 41040 13500 41160
rect 13620 41040 13740 41160
rect 13860 41040 13980 41160
rect 14100 41040 14220 41160
rect 14340 41040 14460 41160
rect 14580 41040 14700 41160
rect 14820 41040 14940 41160
rect 15060 41040 15180 41160
rect 15300 41040 15420 41160
rect 15540 41040 15660 41160
rect 15780 41040 15900 41160
rect 16020 41040 16140 41160
rect 16260 41040 16380 41160
rect 16500 41040 16620 41160
rect 16740 41040 16860 41160
rect 16980 41040 17100 41160
rect 17220 41040 17340 41160
rect 17460 41040 17580 41160
rect 17940 41040 18060 41160
rect 18180 41040 18300 41160
rect 18420 41040 18540 41160
rect 18660 41040 18780 41160
rect 18900 41040 19020 41160
rect 19140 41040 19260 41160
rect 19380 41040 19500 41160
rect 19620 41040 19740 41160
rect 19860 41040 19980 41160
rect 20100 41040 20220 41160
rect 20340 41040 20460 41160
rect 20580 41040 20700 41160
rect 20820 41040 20940 41160
rect 21060 41040 21180 41160
rect 21540 41040 21660 41160
rect 21780 41040 21900 41160
rect 22020 41040 22140 41160
rect 22260 41040 22380 41160
rect 22500 41040 22620 41160
rect 22740 41040 22860 41160
rect 22980 41040 23100 41160
rect 23220 41040 23340 41160
rect 23460 41040 23580 41160
rect 23700 41040 23820 41160
rect 23940 41040 24060 41160
rect 24180 41040 24300 41160
rect 24420 41040 24540 41160
rect 24660 41040 24780 41160
rect 24900 41040 25020 41160
rect 25140 41040 25260 41160
rect 25380 41040 25500 41160
rect 25620 41040 25740 41160
rect 25860 41040 25980 41160
rect 26100 41040 26220 41160
rect 26340 41040 26460 41160
rect 26580 41040 26700 41160
rect 27060 41040 27180 41160
rect 27300 41040 27420 41160
rect 27540 41040 27660 41160
rect 27780 41040 27900 41160
rect 28260 41040 28380 41160
rect 28500 41040 28620 41160
rect 28740 41040 28860 41160
rect 28980 41040 29100 41160
rect 29220 41040 29340 41160
rect 29460 41040 29580 41160
rect 29700 41040 29820 41160
rect 29940 41040 30060 41160
rect 30180 41040 30300 41160
rect 30420 41040 30540 41160
rect 30660 41040 30780 41160
rect 31140 41040 31260 41160
rect 31380 41040 31500 41160
rect 31620 41040 31740 41160
rect 31860 41040 31980 41160
rect 32100 41040 32220 41160
rect 32580 41040 32700 41160
rect 32820 41040 32940 41160
rect 33060 41040 33180 41160
rect 33300 41040 33420 41160
rect 33780 41040 33900 41160
rect 34020 41040 34140 41160
rect 34260 41040 34380 41160
rect 34500 41040 34620 41160
rect 34740 41040 34860 41160
rect 34980 41040 35100 41160
rect 35220 41040 35340 41160
rect 35460 41040 35580 41160
rect 35700 41040 35820 41160
rect 35940 41040 36060 41160
rect 36180 41040 36300 41160
rect 36420 41040 36540 41160
rect 36660 41040 36780 41160
rect 36900 41040 37020 41160
rect 37140 41040 37260 41160
rect 37380 41040 37500 41160
rect 37620 41040 37740 41160
rect 37860 41040 37980 41160
rect 38100 41040 38220 41160
rect 38340 41040 38460 41160
rect 38580 41040 38700 41160
rect 38820 41040 38940 41160
rect 39060 41040 39180 41160
rect 39300 41040 39420 41160
rect 39540 41040 39660 41160
rect 39780 41040 39900 41160
rect 40020 41040 40140 41160
rect 40260 41040 40380 41160
rect 40500 41040 40620 41160
rect 40740 41040 40860 41160
rect 40980 41040 41100 41160
rect 41220 41040 41340 41160
rect 41460 41040 41580 41160
rect 41700 41040 41820 41160
rect 42180 41040 42300 41160
rect 42420 41040 42540 41160
rect 42660 41040 42780 41160
rect 42900 41040 43020 41160
rect 43380 41040 43500 41160
rect 43860 41040 43980 41160
rect 44100 41040 44220 41160
rect 44340 41040 44460 41160
rect 44580 41040 44700 41160
rect 45060 41040 45180 41160
rect 45300 41040 45420 41160
rect 45540 41040 45660 41160
rect 45780 41040 45900 41160
rect 46020 41040 46140 41160
rect 46260 41040 46380 41160
rect 46500 41040 46620 41160
rect 46740 41040 46860 41160
rect 46980 41040 47100 41160
rect 47220 41040 47340 41160
rect 47460 41040 47580 41160
rect 47700 41040 47820 41160
rect 47940 41040 48060 41160
rect 48180 41040 48300 41160
rect 48420 41040 48540 41160
rect 48660 41040 48780 41160
rect 48900 41040 49020 41160
rect 49140 41040 49260 41160
rect 49380 41040 49500 41160
rect 49620 41040 49740 41160
rect 49860 41040 49980 41160
rect 50100 41040 50220 41160
rect 5220 35040 5340 35160
rect 5460 35040 5580 35160
rect 5700 35040 5820 35160
rect 5940 35040 6060 35160
rect 6180 35040 6300 35160
rect 6420 35040 6540 35160
rect 6660 35040 6780 35160
rect 6900 35040 7020 35160
rect 7380 35040 7500 35160
rect 7620 35040 7740 35160
rect 7860 35040 7980 35160
rect 8100 35040 8220 35160
rect 8580 35040 8700 35160
rect 8820 35040 8940 35160
rect 9060 35040 9180 35160
rect 9300 35040 9420 35160
rect 9540 35040 9660 35160
rect 9780 35040 9900 35160
rect 10020 35040 10140 35160
rect 10260 35040 10380 35160
rect 10500 35040 10620 35160
rect 10740 35040 10860 35160
rect 10980 35040 11100 35160
rect 11220 35040 11340 35160
rect 11460 35040 11580 35160
rect 11700 35040 11820 35160
rect 11940 35040 12060 35160
rect 12420 35040 12540 35160
rect 12660 35040 12780 35160
rect 12900 35040 13020 35160
rect 13140 35040 13260 35160
rect 13380 35040 13500 35160
rect 13620 35040 13740 35160
rect 13860 35040 13980 35160
rect 14100 35040 14220 35160
rect 14340 35040 14460 35160
rect 14580 35040 14700 35160
rect 14820 35040 14940 35160
rect 15060 35040 15180 35160
rect 15300 35040 15420 35160
rect 15540 35040 15660 35160
rect 15780 35040 15900 35160
rect 16020 35040 16140 35160
rect 16260 35040 16380 35160
rect 16500 35040 16620 35160
rect 16980 35040 17100 35160
rect 17460 35040 17580 35160
rect 17700 35040 17820 35160
rect 17940 35040 18060 35160
rect 18180 35040 18300 35160
rect 18420 35040 18540 35160
rect 18660 35040 18780 35160
rect 18900 35040 19020 35160
rect 19140 35040 19260 35160
rect 19380 35040 19500 35160
rect 19860 35040 19980 35160
rect 20100 35040 20220 35160
rect 20340 35040 20460 35160
rect 20580 35040 20700 35160
rect 20820 35040 20940 35160
rect 21060 35040 21180 35160
rect 21300 35040 21420 35160
rect 21540 35040 21660 35160
rect 21780 35040 21900 35160
rect 22020 35040 22140 35160
rect 22260 35040 22380 35160
rect 22500 35040 22620 35160
rect 22740 35040 22860 35160
rect 22980 35040 23100 35160
rect 23220 35040 23340 35160
rect 23460 35040 23580 35160
rect 23700 35040 23820 35160
rect 24180 35040 24300 35160
rect 24420 35040 24540 35160
rect 24660 35040 24780 35160
rect 24900 35040 25020 35160
rect 25140 35040 25260 35160
rect 25620 35040 25740 35160
rect 25860 35040 25980 35160
rect 26100 35040 26220 35160
rect 26340 35040 26460 35160
rect 26820 35040 26940 35160
rect 27300 35040 27420 35160
rect 27540 35040 27660 35160
rect 27780 35040 27900 35160
rect 28020 35040 28140 35160
rect 28260 35040 28380 35160
rect 28500 35040 28620 35160
rect 28740 35040 28860 35160
rect 28980 35040 29100 35160
rect 29220 35040 29340 35160
rect 29460 35040 29580 35160
rect 29700 35040 29820 35160
rect 29940 35040 30060 35160
rect 30180 35040 30300 35160
rect 30420 35040 30540 35160
rect 30660 35040 30780 35160
rect 30900 35040 31020 35160
rect 31140 35040 31260 35160
rect 31620 35040 31740 35160
rect 31860 35040 31980 35160
rect 32340 35040 32460 35160
rect 32820 35040 32940 35160
rect 33060 35040 33180 35160
rect 33300 35040 33420 35160
rect 33540 35040 33660 35160
rect 33780 35040 33900 35160
rect 34020 35040 34140 35160
rect 34260 35040 34380 35160
rect 34500 35040 34620 35160
rect 34980 35040 35100 35160
rect 35220 35040 35340 35160
rect 35460 35040 35580 35160
rect 35700 35040 35820 35160
rect 35940 35040 36060 35160
rect 36180 35040 36300 35160
rect 36420 35040 36540 35160
rect 36660 35040 36780 35160
rect 36900 35040 37020 35160
rect 37140 35040 37260 35160
rect 37380 35040 37500 35160
rect 37620 35040 37740 35160
rect 37860 35040 37980 35160
rect 38100 35040 38220 35160
rect 38340 35040 38460 35160
rect 38580 35040 38700 35160
rect 38820 35040 38940 35160
rect 39300 35040 39420 35160
rect 39540 35040 39660 35160
rect 39780 35040 39900 35160
rect 40020 35040 40140 35160
rect 40500 35040 40620 35160
rect 40980 35040 41100 35160
rect 41220 35040 41340 35160
rect 41460 35040 41580 35160
rect 41940 35040 42060 35160
rect 42180 35040 42300 35160
rect 42420 35040 42540 35160
rect 42660 35040 42780 35160
rect 42900 35040 43020 35160
rect 43140 35040 43260 35160
rect 43380 35040 43500 35160
rect 43860 35040 43980 35160
rect 44100 35040 44220 35160
rect 44340 35040 44460 35160
rect 44580 35040 44700 35160
rect 44820 35040 44940 35160
rect 45060 35040 45180 35160
rect 45300 35040 45420 35160
rect 45540 35040 45660 35160
rect 45780 35040 45900 35160
rect 46020 35040 46140 35160
rect 46500 35040 46620 35160
rect 46740 35040 46860 35160
rect 46980 35040 47100 35160
rect 47220 35040 47340 35160
rect 47460 35040 47580 35160
rect 47700 35040 47820 35160
rect 47940 35040 48060 35160
rect 48180 35040 48300 35160
rect 48420 35040 48540 35160
rect 48660 35040 48780 35160
rect 48900 35040 49020 35160
rect 49140 35040 49260 35160
rect 49380 35040 49500 35160
rect 49620 35040 49740 35160
rect 49860 35040 49980 35160
rect 50100 35040 50220 35160
rect 5220 29040 5340 29160
rect 5460 29040 5580 29160
rect 5700 29040 5820 29160
rect 5940 29040 6060 29160
rect 6180 29040 6300 29160
rect 6420 29040 6540 29160
rect 6660 29040 6780 29160
rect 6900 29040 7020 29160
rect 7140 29040 7260 29160
rect 7380 29040 7500 29160
rect 7620 29040 7740 29160
rect 7860 29040 7980 29160
rect 8340 29040 8460 29160
rect 8580 29040 8700 29160
rect 8820 29040 8940 29160
rect 9060 29040 9180 29160
rect 9300 29040 9420 29160
rect 9540 29040 9660 29160
rect 9780 29040 9900 29160
rect 10020 29040 10140 29160
rect 10260 29040 10380 29160
rect 10500 29040 10620 29160
rect 10740 29040 10860 29160
rect 10980 29040 11100 29160
rect 11460 29040 11580 29160
rect 11940 29040 12060 29160
rect 12420 29040 12540 29160
rect 12660 29040 12780 29160
rect 12900 29040 13020 29160
rect 13140 29040 13260 29160
rect 13380 29040 13500 29160
rect 13620 29040 13740 29160
rect 13860 29040 13980 29160
rect 14100 29040 14220 29160
rect 14340 29040 14460 29160
rect 14580 29040 14700 29160
rect 14820 29040 14940 29160
rect 15060 29040 15180 29160
rect 15300 29040 15420 29160
rect 15540 29040 15660 29160
rect 15780 29040 15900 29160
rect 16020 29040 16140 29160
rect 16260 29040 16380 29160
rect 16500 29040 16620 29160
rect 16740 29040 16860 29160
rect 16980 29040 17100 29160
rect 17220 29040 17340 29160
rect 17460 29040 17580 29160
rect 17700 29040 17820 29160
rect 17940 29040 18060 29160
rect 18420 29040 18540 29160
rect 18660 29040 18780 29160
rect 18900 29040 19020 29160
rect 19140 29040 19260 29160
rect 19620 29040 19740 29160
rect 20100 29040 20220 29160
rect 20340 29040 20460 29160
rect 20580 29040 20700 29160
rect 20820 29040 20940 29160
rect 21060 29040 21180 29160
rect 21300 29040 21420 29160
rect 21540 29040 21660 29160
rect 21780 29040 21900 29160
rect 22020 29040 22140 29160
rect 22500 29040 22620 29160
rect 22740 29040 22860 29160
rect 22980 29040 23100 29160
rect 23220 29040 23340 29160
rect 23460 29040 23580 29160
rect 23700 29040 23820 29160
rect 23940 29040 24060 29160
rect 24180 29040 24300 29160
rect 24420 29040 24540 29160
rect 24660 29040 24780 29160
rect 24900 29040 25020 29160
rect 25140 29040 25260 29160
rect 25380 29040 25500 29160
rect 25620 29040 25740 29160
rect 25860 29040 25980 29160
rect 26100 29040 26220 29160
rect 26340 29040 26460 29160
rect 26820 29040 26940 29160
rect 27060 29040 27180 29160
rect 27300 29040 27420 29160
rect 27540 29040 27660 29160
rect 27780 29040 27900 29160
rect 28020 29040 28140 29160
rect 28260 29040 28380 29160
rect 28500 29040 28620 29160
rect 28740 29040 28860 29160
rect 29220 29040 29340 29160
rect 29460 29040 29580 29160
rect 29700 29040 29820 29160
rect 29940 29040 30060 29160
rect 30180 29040 30300 29160
rect 30420 29040 30540 29160
rect 30660 29040 30780 29160
rect 30900 29040 31020 29160
rect 31140 29040 31260 29160
rect 31380 29040 31500 29160
rect 31620 29040 31740 29160
rect 31860 29040 31980 29160
rect 32100 29040 32220 29160
rect 32340 29040 32460 29160
rect 32580 29040 32700 29160
rect 32820 29040 32940 29160
rect 33060 29040 33180 29160
rect 33300 29040 33420 29160
rect 33540 29040 33660 29160
rect 33780 29040 33900 29160
rect 34020 29040 34140 29160
rect 34260 29040 34380 29160
rect 34500 29040 34620 29160
rect 34740 29040 34860 29160
rect 34980 29040 35100 29160
rect 35220 29040 35340 29160
rect 35460 29040 35580 29160
rect 35700 29040 35820 29160
rect 35940 29040 36060 29160
rect 36420 29040 36540 29160
rect 36660 29040 36780 29160
rect 36900 29040 37020 29160
rect 37140 29040 37260 29160
rect 37380 29040 37500 29160
rect 37620 29040 37740 29160
rect 38100 29040 38220 29160
rect 38340 29040 38460 29160
rect 38580 29040 38700 29160
rect 38820 29040 38940 29160
rect 39060 29040 39180 29160
rect 39300 29040 39420 29160
rect 39540 29040 39660 29160
rect 39780 29040 39900 29160
rect 40020 29040 40140 29160
rect 40260 29040 40380 29160
rect 40500 29040 40620 29160
rect 40980 29040 41100 29160
rect 41220 29040 41340 29160
rect 41460 29040 41580 29160
rect 41700 29040 41820 29160
rect 41940 29040 42060 29160
rect 42180 29040 42300 29160
rect 42420 29040 42540 29160
rect 42660 29040 42780 29160
rect 42900 29040 43020 29160
rect 43380 29040 43500 29160
rect 43860 29040 43980 29160
rect 44100 29040 44220 29160
rect 44340 29040 44460 29160
rect 44820 29040 44940 29160
rect 45300 29040 45420 29160
rect 45540 29040 45660 29160
rect 45780 29040 45900 29160
rect 46020 29040 46140 29160
rect 46260 29040 46380 29160
rect 46740 29040 46860 29160
rect 46980 29040 47100 29160
rect 47220 29040 47340 29160
rect 47460 29040 47580 29160
rect 47700 29040 47820 29160
rect 47940 29040 48060 29160
rect 48420 29040 48540 29160
rect 48900 29040 49020 29160
rect 49140 29040 49260 29160
rect 49380 29040 49500 29160
rect 49620 29040 49740 29160
rect 49860 29040 49980 29160
rect 50100 29040 50220 29160
rect 5220 23040 5340 23160
rect 5700 23040 5820 23160
rect 6180 23040 6300 23160
rect 6660 23040 6780 23160
rect 6900 23040 7020 23160
rect 7140 23040 7260 23160
rect 7380 23040 7500 23160
rect 7620 23040 7740 23160
rect 7860 23040 7980 23160
rect 8100 23040 8220 23160
rect 8580 23040 8700 23160
rect 8820 23040 8940 23160
rect 9060 23040 9180 23160
rect 9300 23040 9420 23160
rect 9540 23040 9660 23160
rect 9780 23040 9900 23160
rect 10020 23040 10140 23160
rect 10260 23040 10380 23160
rect 10500 23040 10620 23160
rect 10740 23040 10860 23160
rect 10980 23040 11100 23160
rect 11220 23040 11340 23160
rect 11460 23040 11580 23160
rect 11700 23040 11820 23160
rect 11940 23040 12060 23160
rect 12180 23040 12300 23160
rect 12420 23040 12540 23160
rect 12660 23040 12780 23160
rect 12900 23040 13020 23160
rect 13140 23040 13260 23160
rect 13380 23040 13500 23160
rect 13620 23040 13740 23160
rect 13860 23040 13980 23160
rect 14100 23040 14220 23160
rect 14340 23040 14460 23160
rect 14580 23040 14700 23160
rect 14820 23040 14940 23160
rect 15060 23040 15180 23160
rect 15300 23040 15420 23160
rect 15540 23040 15660 23160
rect 15780 23040 15900 23160
rect 16020 23040 16140 23160
rect 16260 23040 16380 23160
rect 16500 23040 16620 23160
rect 16740 23040 16860 23160
rect 16980 23040 17100 23160
rect 17220 23040 17340 23160
rect 17460 23040 17580 23160
rect 17700 23040 17820 23160
rect 17940 23040 18060 23160
rect 18180 23040 18300 23160
rect 18420 23040 18540 23160
rect 18660 23040 18780 23160
rect 18900 23040 19020 23160
rect 19140 23040 19260 23160
rect 19380 23040 19500 23160
rect 19620 23040 19740 23160
rect 19860 23040 19980 23160
rect 20100 23040 20220 23160
rect 20340 23040 20460 23160
rect 20580 23040 20700 23160
rect 20820 23040 20940 23160
rect 21060 23040 21180 23160
rect 21300 23040 21420 23160
rect 21540 23040 21660 23160
rect 21780 23040 21900 23160
rect 22020 23040 22140 23160
rect 22260 23040 22380 23160
rect 22500 23040 22620 23160
rect 22740 23040 22860 23160
rect 22980 23040 23100 23160
rect 23220 23040 23340 23160
rect 23460 23040 23580 23160
rect 23700 23040 23820 23160
rect 23940 23040 24060 23160
rect 24180 23040 24300 23160
rect 24420 23040 24540 23160
rect 24660 23040 24780 23160
rect 24900 23040 25020 23160
rect 25140 23040 25260 23160
rect 25380 23040 25500 23160
rect 25620 23040 25740 23160
rect 25860 23040 25980 23160
rect 26100 23040 26220 23160
rect 26580 23040 26700 23160
rect 27060 23040 27180 23160
rect 27300 23040 27420 23160
rect 27540 23040 27660 23160
rect 27780 23040 27900 23160
rect 28260 23040 28380 23160
rect 28740 23040 28860 23160
rect 28980 23040 29100 23160
rect 29220 23040 29340 23160
rect 29460 23040 29580 23160
rect 29700 23040 29820 23160
rect 29940 23040 30060 23160
rect 30180 23040 30300 23160
rect 30660 23040 30780 23160
rect 30900 23040 31020 23160
rect 31140 23040 31260 23160
rect 31380 23040 31500 23160
rect 31620 23040 31740 23160
rect 31860 23040 31980 23160
rect 32100 23040 32220 23160
rect 32340 23040 32460 23160
rect 32580 23040 32700 23160
rect 32820 23040 32940 23160
rect 33060 23040 33180 23160
rect 33540 23040 33660 23160
rect 33780 23040 33900 23160
rect 34020 23040 34140 23160
rect 34260 23040 34380 23160
rect 34500 23040 34620 23160
rect 34980 23040 35100 23160
rect 35220 23040 35340 23160
rect 35460 23040 35580 23160
rect 35700 23040 35820 23160
rect 35940 23040 36060 23160
rect 36180 23040 36300 23160
rect 36420 23040 36540 23160
rect 36660 23040 36780 23160
rect 36900 23040 37020 23160
rect 37140 23040 37260 23160
rect 37380 23040 37500 23160
rect 37620 23040 37740 23160
rect 37860 23040 37980 23160
rect 38100 23040 38220 23160
rect 38340 23040 38460 23160
rect 38580 23040 38700 23160
rect 38820 23040 38940 23160
rect 39300 23040 39420 23160
rect 39540 23040 39660 23160
rect 39780 23040 39900 23160
rect 40020 23040 40140 23160
rect 40260 23040 40380 23160
rect 40740 23040 40860 23160
rect 40980 23040 41100 23160
rect 41220 23040 41340 23160
rect 41460 23040 41580 23160
rect 41700 23040 41820 23160
rect 41940 23040 42060 23160
rect 42180 23040 42300 23160
rect 42420 23040 42540 23160
rect 42660 23040 42780 23160
rect 42900 23040 43020 23160
rect 43140 23040 43260 23160
rect 43620 23040 43740 23160
rect 43860 23040 43980 23160
rect 44100 23040 44220 23160
rect 44340 23040 44460 23160
rect 44580 23040 44700 23160
rect 44820 23040 44940 23160
rect 45060 23040 45180 23160
rect 45300 23040 45420 23160
rect 45540 23040 45660 23160
rect 45780 23040 45900 23160
rect 46020 23040 46140 23160
rect 46260 23040 46380 23160
rect 46500 23040 46620 23160
rect 46740 23040 46860 23160
rect 46980 23040 47100 23160
rect 47220 23040 47340 23160
rect 47460 23040 47580 23160
rect 47700 23040 47820 23160
rect 47940 23040 48060 23160
rect 48180 23040 48300 23160
rect 48420 23040 48540 23160
rect 48660 23040 48780 23160
rect 48900 23040 49020 23160
rect 49140 23040 49260 23160
rect 49380 23040 49500 23160
rect 49620 23040 49740 23160
rect 49860 23040 49980 23160
rect 50100 23040 50220 23160
rect 5220 17040 5340 17160
rect 5460 17040 5580 17160
rect 5700 17040 5820 17160
rect 5940 17040 6060 17160
rect 6180 17040 6300 17160
rect 6420 17040 6540 17160
rect 6660 17040 6780 17160
rect 6900 17040 7020 17160
rect 7140 17040 7260 17160
rect 7380 17040 7500 17160
rect 7620 17040 7740 17160
rect 7860 17040 7980 17160
rect 8100 17040 8220 17160
rect 8340 17040 8460 17160
rect 8580 17040 8700 17160
rect 8820 17040 8940 17160
rect 9060 17040 9180 17160
rect 9300 17040 9420 17160
rect 9540 17040 9660 17160
rect 9780 17040 9900 17160
rect 10020 17040 10140 17160
rect 10260 17040 10380 17160
rect 10500 17040 10620 17160
rect 10740 17040 10860 17160
rect 10980 17040 11100 17160
rect 11220 17040 11340 17160
rect 11460 17040 11580 17160
rect 11940 17040 12060 17160
rect 12420 17040 12540 17160
rect 12660 17040 12780 17160
rect 12900 17040 13020 17160
rect 13140 17040 13260 17160
rect 13380 17040 13500 17160
rect 13620 17040 13740 17160
rect 13860 17040 13980 17160
rect 14100 17040 14220 17160
rect 14340 17040 14460 17160
rect 14580 17040 14700 17160
rect 14820 17040 14940 17160
rect 15060 17040 15180 17160
rect 15300 17040 15420 17160
rect 15780 17040 15900 17160
rect 16260 17040 16380 17160
rect 16500 17040 16620 17160
rect 16740 17040 16860 17160
rect 16980 17040 17100 17160
rect 17220 17040 17340 17160
rect 17460 17040 17580 17160
rect 17700 17040 17820 17160
rect 17940 17040 18060 17160
rect 18180 17040 18300 17160
rect 18420 17040 18540 17160
rect 18660 17040 18780 17160
rect 18900 17040 19020 17160
rect 19140 17040 19260 17160
rect 19380 17040 19500 17160
rect 19620 17040 19740 17160
rect 19860 17040 19980 17160
rect 20100 17040 20220 17160
rect 20340 17040 20460 17160
rect 20580 17040 20700 17160
rect 20820 17040 20940 17160
rect 21060 17040 21180 17160
rect 21300 17040 21420 17160
rect 21540 17040 21660 17160
rect 21780 17040 21900 17160
rect 22020 17040 22140 17160
rect 22500 17040 22620 17160
rect 22740 17040 22860 17160
rect 22980 17040 23100 17160
rect 23220 17040 23340 17160
rect 23460 17040 23580 17160
rect 23940 17040 24060 17160
rect 24180 17040 24300 17160
rect 24420 17040 24540 17160
rect 24660 17040 24780 17160
rect 24900 17040 25020 17160
rect 25380 17040 25500 17160
rect 25620 17040 25740 17160
rect 25860 17040 25980 17160
rect 26100 17040 26220 17160
rect 26340 17040 26460 17160
rect 26580 17040 26700 17160
rect 26820 17040 26940 17160
rect 27300 17040 27420 17160
rect 27540 17040 27660 17160
rect 27780 17040 27900 17160
rect 28020 17040 28140 17160
rect 28260 17040 28380 17160
rect 28500 17040 28620 17160
rect 28740 17040 28860 17160
rect 28980 17040 29100 17160
rect 29220 17040 29340 17160
rect 29460 17040 29580 17160
rect 29700 17040 29820 17160
rect 29940 17040 30060 17160
rect 30180 17040 30300 17160
rect 30420 17040 30540 17160
rect 30900 17040 31020 17160
rect 31140 17040 31260 17160
rect 31380 17040 31500 17160
rect 31620 17040 31740 17160
rect 31860 17040 31980 17160
rect 32100 17040 32220 17160
rect 32340 17040 32460 17160
rect 32580 17040 32700 17160
rect 32820 17040 32940 17160
rect 33060 17040 33180 17160
rect 33540 17040 33660 17160
rect 33780 17040 33900 17160
rect 34020 17040 34140 17160
rect 34260 17040 34380 17160
rect 34500 17040 34620 17160
rect 34740 17040 34860 17160
rect 34980 17040 35100 17160
rect 35220 17040 35340 17160
rect 35460 17040 35580 17160
rect 35700 17040 35820 17160
rect 35940 17040 36060 17160
rect 36180 17040 36300 17160
rect 36420 17040 36540 17160
rect 36660 17040 36780 17160
rect 36900 17040 37020 17160
rect 37140 17040 37260 17160
rect 37380 17040 37500 17160
rect 37620 17040 37740 17160
rect 37860 17040 37980 17160
rect 38100 17040 38220 17160
rect 38340 17040 38460 17160
rect 38580 17040 38700 17160
rect 38820 17040 38940 17160
rect 39300 17040 39420 17160
rect 39540 17040 39660 17160
rect 39780 17040 39900 17160
rect 40020 17040 40140 17160
rect 40260 17040 40380 17160
rect 40500 17040 40620 17160
rect 40740 17040 40860 17160
rect 40980 17040 41100 17160
rect 41220 17040 41340 17160
rect 41460 17040 41580 17160
rect 41940 17040 42060 17160
rect 42180 17040 42300 17160
rect 42420 17040 42540 17160
rect 42660 17040 42780 17160
rect 42900 17040 43020 17160
rect 43140 17040 43260 17160
rect 43380 17040 43500 17160
rect 43620 17040 43740 17160
rect 43860 17040 43980 17160
rect 44100 17040 44220 17160
rect 44340 17040 44460 17160
rect 44820 17040 44940 17160
rect 45300 17040 45420 17160
rect 45540 17040 45660 17160
rect 45780 17040 45900 17160
rect 46020 17040 46140 17160
rect 46500 17040 46620 17160
rect 46740 17040 46860 17160
rect 46980 17040 47100 17160
rect 47220 17040 47340 17160
rect 47460 17040 47580 17160
rect 47700 17040 47820 17160
rect 47940 17040 48060 17160
rect 48180 17040 48300 17160
rect 48420 17040 48540 17160
rect 48660 17040 48780 17160
rect 48900 17040 49020 17160
rect 49380 17040 49500 17160
rect 49860 17040 49980 17160
rect 50100 17040 50220 17160
rect 5220 11040 5340 11160
rect 5460 11040 5580 11160
rect 5700 11040 5820 11160
rect 5940 11040 6060 11160
rect 6180 11040 6300 11160
rect 6420 11040 6540 11160
rect 6660 11040 6780 11160
rect 6900 11040 7020 11160
rect 7140 11040 7260 11160
rect 7380 11040 7500 11160
rect 7620 11040 7740 11160
rect 7860 11040 7980 11160
rect 8100 11040 8220 11160
rect 8340 11040 8460 11160
rect 8580 11040 8700 11160
rect 8820 11040 8940 11160
rect 9060 11040 9180 11160
rect 9300 11040 9420 11160
rect 9540 11040 9660 11160
rect 9780 11040 9900 11160
rect 10020 11040 10140 11160
rect 10260 11040 10380 11160
rect 10500 11040 10620 11160
rect 10740 11040 10860 11160
rect 10980 11040 11100 11160
rect 11220 11040 11340 11160
rect 11460 11040 11580 11160
rect 11700 11040 11820 11160
rect 11940 11040 12060 11160
rect 12180 11040 12300 11160
rect 12420 11040 12540 11160
rect 12660 11040 12780 11160
rect 12900 11040 13020 11160
rect 13140 11040 13260 11160
rect 13380 11040 13500 11160
rect 13620 11040 13740 11160
rect 13860 11040 13980 11160
rect 14100 11040 14220 11160
rect 14340 11040 14460 11160
rect 14580 11040 14700 11160
rect 14820 11040 14940 11160
rect 15060 11040 15180 11160
rect 15300 11040 15420 11160
rect 15540 11040 15660 11160
rect 15780 11040 15900 11160
rect 16020 11040 16140 11160
rect 16260 11040 16380 11160
rect 16740 11040 16860 11160
rect 16980 11040 17100 11160
rect 17220 11040 17340 11160
rect 17460 11040 17580 11160
rect 17700 11040 17820 11160
rect 17940 11040 18060 11160
rect 18180 11040 18300 11160
rect 18420 11040 18540 11160
rect 18660 11040 18780 11160
rect 18900 11040 19020 11160
rect 19140 11040 19260 11160
rect 19380 11040 19500 11160
rect 19860 11040 19980 11160
rect 20340 11040 20460 11160
rect 20820 11040 20940 11160
rect 21060 11040 21180 11160
rect 21300 11040 21420 11160
rect 21540 11040 21660 11160
rect 21780 11040 21900 11160
rect 22020 11040 22140 11160
rect 22260 11040 22380 11160
rect 22500 11040 22620 11160
rect 22740 11040 22860 11160
rect 22980 11040 23100 11160
rect 23220 11040 23340 11160
rect 23460 11040 23580 11160
rect 23700 11040 23820 11160
rect 23940 11040 24060 11160
rect 24180 11040 24300 11160
rect 24420 11040 24540 11160
rect 24660 11040 24780 11160
rect 24900 11040 25020 11160
rect 25140 11040 25260 11160
rect 25380 11040 25500 11160
rect 25860 11040 25980 11160
rect 26100 11040 26220 11160
rect 26340 11040 26460 11160
rect 26580 11040 26700 11160
rect 26820 11040 26940 11160
rect 27060 11040 27180 11160
rect 27300 11040 27420 11160
rect 27540 11040 27660 11160
rect 27780 11040 27900 11160
rect 28020 11040 28140 11160
rect 28260 11040 28380 11160
rect 28500 11040 28620 11160
rect 28740 11040 28860 11160
rect 28980 11040 29100 11160
rect 29220 11040 29340 11160
rect 29460 11040 29580 11160
rect 29700 11040 29820 11160
rect 29940 11040 30060 11160
rect 30180 11040 30300 11160
rect 30420 11040 30540 11160
rect 30660 11040 30780 11160
rect 30900 11040 31020 11160
rect 31140 11040 31260 11160
rect 31380 11040 31500 11160
rect 31620 11040 31740 11160
rect 31860 11040 31980 11160
rect 32100 11040 32220 11160
rect 32580 11040 32700 11160
rect 32820 11040 32940 11160
rect 33060 11040 33180 11160
rect 33300 11040 33420 11160
rect 33780 11040 33900 11160
rect 34260 11040 34380 11160
rect 34500 11040 34620 11160
rect 34740 11040 34860 11160
rect 34980 11040 35100 11160
rect 35220 11040 35340 11160
rect 35460 11040 35580 11160
rect 35700 11040 35820 11160
rect 35940 11040 36060 11160
rect 36420 11040 36540 11160
rect 36660 11040 36780 11160
rect 36900 11040 37020 11160
rect 37140 11040 37260 11160
rect 37380 11040 37500 11160
rect 37620 11040 37740 11160
rect 37860 11040 37980 11160
rect 38100 11040 38220 11160
rect 38340 11040 38460 11160
rect 38580 11040 38700 11160
rect 38820 11040 38940 11160
rect 39300 11040 39420 11160
rect 39540 11040 39660 11160
rect 39780 11040 39900 11160
rect 40020 11040 40140 11160
rect 40260 11040 40380 11160
rect 40500 11040 40620 11160
rect 40740 11040 40860 11160
rect 40980 11040 41100 11160
rect 41220 11040 41340 11160
rect 41460 11040 41580 11160
rect 41940 11040 42060 11160
rect 42180 11040 42300 11160
rect 42420 11040 42540 11160
rect 42660 11040 42780 11160
rect 42900 11040 43020 11160
rect 43140 11040 43260 11160
rect 43380 11040 43500 11160
rect 43620 11040 43740 11160
rect 43860 11040 43980 11160
rect 44100 11040 44220 11160
rect 44340 11040 44460 11160
rect 44580 11040 44700 11160
rect 44820 11040 44940 11160
rect 45060 11040 45180 11160
rect 45300 11040 45420 11160
rect 45540 11040 45660 11160
rect 45780 11040 45900 11160
rect 46020 11040 46140 11160
rect 46500 11040 46620 11160
rect 46740 11040 46860 11160
rect 46980 11040 47100 11160
rect 47220 11040 47340 11160
rect 47460 11040 47580 11160
rect 47700 11040 47820 11160
rect 47940 11040 48060 11160
rect 48180 11040 48300 11160
rect 48420 11040 48540 11160
rect 48660 11040 48780 11160
rect 48900 11040 49020 11160
rect 49140 11040 49260 11160
rect 49380 11040 49500 11160
rect 49620 11040 49740 11160
rect 49860 11040 49980 11160
rect 50100 11040 50220 11160
rect 5220 5040 5340 5160
rect 5460 5040 5580 5160
rect 5700 5040 5820 5160
rect 6180 5040 6300 5160
rect 6660 5040 6780 5160
rect 7140 5040 7260 5160
rect 7380 5040 7500 5160
rect 7620 5040 7740 5160
rect 7860 5040 7980 5160
rect 8340 5040 8460 5160
rect 8580 5040 8700 5160
rect 9060 5040 9180 5160
rect 9540 5040 9660 5160
rect 9780 5040 9900 5160
rect 10260 5040 10380 5160
rect 10500 5040 10620 5160
rect 10740 5040 10860 5160
rect 11220 5040 11340 5160
rect 11700 5040 11820 5160
rect 11940 5040 12060 5160
rect 12180 5040 12300 5160
rect 12660 5040 12780 5160
rect 12900 5040 13020 5160
rect 13140 5040 13260 5160
rect 13380 5040 13500 5160
rect 13620 5040 13740 5160
rect 14100 5040 14220 5160
rect 14580 5040 14700 5160
rect 14820 5040 14940 5160
rect 15060 5040 15180 5160
rect 15300 5040 15420 5160
rect 15780 5040 15900 5160
rect 16020 5040 16140 5160
rect 16260 5040 16380 5160
rect 16500 5040 16620 5160
rect 16740 5040 16860 5160
rect 16980 5040 17100 5160
rect 17220 5040 17340 5160
rect 17460 5040 17580 5160
rect 17700 5040 17820 5160
rect 17940 5040 18060 5160
rect 18420 5040 18540 5160
rect 18660 5040 18780 5160
rect 18900 5040 19020 5160
rect 19140 5040 19260 5160
rect 19380 5040 19500 5160
rect 19620 5040 19740 5160
rect 19860 5040 19980 5160
rect 20100 5040 20220 5160
rect 20340 5040 20460 5160
rect 20580 5040 20700 5160
rect 21060 5040 21180 5160
rect 21300 5040 21420 5160
rect 21540 5040 21660 5160
rect 21780 5040 21900 5160
rect 22020 5040 22140 5160
rect 22260 5040 22380 5160
rect 22500 5040 22620 5160
rect 22740 5040 22860 5160
rect 22980 5040 23100 5160
rect 23220 5040 23340 5160
rect 23700 5040 23820 5160
rect 23940 5040 24060 5160
rect 24180 5040 24300 5160
rect 24420 5040 24540 5160
rect 24660 5040 24780 5160
rect 24900 5040 25020 5160
rect 25140 5040 25260 5160
rect 25380 5040 25500 5160
rect 25620 5040 25740 5160
rect 26100 5040 26220 5160
rect 26580 5040 26700 5160
rect 27060 5040 27180 5160
rect 27300 5040 27420 5160
rect 27540 5040 27660 5160
rect 27780 5040 27900 5160
rect 28260 5040 28380 5160
rect 28500 5040 28620 5160
rect 28740 5040 28860 5160
rect 28980 5040 29100 5160
rect 29460 5040 29580 5160
rect 29700 5040 29820 5160
rect 29940 5040 30060 5160
rect 30420 5040 30540 5160
rect 30900 5040 31020 5160
rect 31380 5040 31500 5160
rect 31620 5040 31740 5160
rect 31860 5040 31980 5160
rect 32340 5040 32460 5160
rect 32820 5040 32940 5160
rect 33060 5040 33180 5160
rect 33540 5040 33660 5160
rect 33780 5040 33900 5160
rect 34020 5040 34140 5160
rect 34260 5040 34380 5160
rect 34500 5040 34620 5160
rect 34740 5040 34860 5160
rect 35220 5040 35340 5160
rect 35460 5040 35580 5160
rect 35700 5040 35820 5160
rect 35940 5040 36060 5160
rect 36420 5040 36540 5160
rect 36660 5040 36780 5160
rect 36900 5040 37020 5160
rect 37140 5040 37260 5160
rect 37380 5040 37500 5160
rect 37860 5040 37980 5160
rect 38340 5040 38460 5160
rect 38580 5040 38700 5160
rect 38820 5040 38940 5160
rect 39300 5040 39420 5160
rect 39540 5040 39660 5160
rect 39780 5040 39900 5160
rect 40020 5040 40140 5160
rect 40260 5040 40380 5160
rect 40740 5040 40860 5160
rect 40980 5040 41100 5160
rect 41220 5040 41340 5160
rect 41460 5040 41580 5160
rect 41700 5040 41820 5160
rect 41940 5040 42060 5160
rect 42180 5040 42300 5160
rect 42420 5040 42540 5160
rect 42660 5040 42780 5160
rect 42900 5040 43020 5160
rect 43140 5040 43260 5160
rect 43620 5040 43740 5160
rect 43860 5040 43980 5160
rect 44100 5040 44220 5160
rect 44340 5040 44460 5160
rect 44820 5040 44940 5160
rect 45300 5040 45420 5160
rect 45540 5040 45660 5160
rect 45780 5040 45900 5160
rect 46020 5040 46140 5160
rect 46260 5040 46380 5160
rect 46740 5040 46860 5160
rect 46980 5040 47100 5160
rect 47220 5040 47340 5160
rect 47700 5040 47820 5160
rect 48180 5040 48300 5160
rect 48420 5040 48540 5160
rect 48660 5040 48780 5160
rect 48900 5040 49020 5160
rect 49140 5040 49260 5160
rect 49380 5040 49500 5160
rect 49620 5040 49740 5160
rect 49860 5040 49980 5160
rect 50100 5040 50220 5160
<< polysilicon >>
rect 5730 43920 5790 43980
rect 5970 43920 6030 43980
rect 6210 43920 6270 43980
rect 6930 43920 6990 43980
rect 7080 43920 7140 43980
rect 7890 43920 7950 43980
rect 8130 43920 8190 43980
rect 8370 43920 8430 43980
rect 9090 43920 9150 43980
rect 9360 43920 9420 43980
rect 9510 43920 9570 43980
rect 9870 43920 9930 43980
rect 10020 43920 10080 43980
rect 10290 43920 10350 43980
rect 11010 43920 11070 43980
rect 11250 43920 11310 43980
rect 12450 43920 12510 43980
rect 12690 43920 12750 43980
rect 13890 43920 13950 43980
rect 14130 43920 14190 43980
rect 14370 43920 14430 43980
rect 15570 43920 15630 43980
rect 15720 43920 15780 43980
rect 17250 43920 17310 43980
rect 17490 43920 17550 43980
rect 17730 43920 17790 43980
rect 19410 43920 19470 43980
rect 19680 43920 19740 43980
rect 19830 43920 19890 43980
rect 20190 43920 20250 43980
rect 20340 43920 20400 43980
rect 20610 43920 20670 43980
rect 21330 43920 21390 43980
rect 22770 43920 22830 43980
rect 23040 43920 23100 43980
rect 23190 43920 23250 43980
rect 23550 43920 23610 43980
rect 23700 43920 23760 43980
rect 23970 43920 24030 43980
rect 25170 43920 25230 43980
rect 25410 43920 25470 43980
rect 25650 43920 25710 43980
rect 26850 43920 26910 43980
rect 27000 43920 27060 43980
rect 28050 43920 28110 43980
rect 28290 43920 28350 43980
rect 28530 43920 28590 43980
rect 29250 43920 29310 43980
rect 29400 43920 29460 43980
rect 30450 43920 30510 43980
rect 30690 43920 30750 43980
rect 30930 43920 30990 43980
rect 31890 43920 31950 43980
rect 32130 43920 32190 43980
rect 32370 43920 32430 43980
rect 33420 43920 33480 43980
rect 33570 43920 33630 43980
rect 34770 43920 34830 43980
rect 35010 43920 35070 43980
rect 35970 43920 36030 43980
rect 36240 43920 36300 43980
rect 36390 43920 36450 43980
rect 36750 43920 36810 43980
rect 36900 43920 36960 43980
rect 37170 43920 37230 43980
rect 37890 43920 37950 43980
rect 38130 43920 38190 43980
rect 38370 43920 38430 43980
rect 39570 43920 39630 43980
rect 39840 43920 39900 43980
rect 39990 43920 40050 43980
rect 40350 43920 40410 43980
rect 40500 43920 40560 43980
rect 40770 43920 40830 43980
rect 41970 43920 42030 43980
rect 43170 43920 43230 43980
rect 43410 43920 43470 43980
rect 43650 43920 43710 43980
rect 44370 43920 44430 43980
rect 44610 43920 44670 43980
rect 44850 43920 44910 43980
rect 45330 43920 45390 43980
rect 45810 43920 45870 43980
rect 46080 43920 46140 43980
rect 46230 43920 46290 43980
rect 46590 43920 46650 43980
rect 46740 43920 46800 43980
rect 47010 43920 47070 43980
rect 47490 43920 47550 43980
rect 47760 43920 47820 43980
rect 47910 43920 47970 43980
rect 48270 43920 48330 43980
rect 48420 43920 48480 43980
rect 48690 43920 48750 43980
rect 5730 42210 5790 43320
rect 5970 42930 6030 43320
rect 6210 43170 6270 43320
rect 6930 43230 6990 43320
rect 7080 43290 7140 43320
rect 7080 43230 7230 43290
rect 6900 43110 6990 43230
rect 5970 42810 6060 42930
rect 5970 42570 6030 42810
rect 6300 42690 6360 43110
rect 6210 42630 6360 42690
rect 5970 42510 6120 42570
rect 6060 42480 6120 42510
rect 6210 42480 6270 42630
rect 5820 41880 5880 42150
rect 6930 41880 6990 43110
rect 7170 42390 7230 43230
rect 7170 42270 7260 42390
rect 7170 41880 7230 42270
rect 7890 42210 7950 43320
rect 8130 42930 8190 43320
rect 8370 43170 8430 43320
rect 9090 43110 9150 43320
rect 9360 43290 9420 43320
rect 9300 43230 9420 43290
rect 9510 43290 9570 43320
rect 9870 43290 9930 43320
rect 8130 42810 8220 42930
rect 8130 42570 8190 42810
rect 8460 42690 8520 43110
rect 8370 42630 8520 42690
rect 8130 42510 8280 42570
rect 8220 42480 8280 42510
rect 8370 42480 8430 42630
rect 9090 42480 9150 42990
rect 9300 42810 9360 43230
rect 9510 43170 9540 43290
rect 9780 43230 9930 43290
rect 10020 43290 10080 43320
rect 10290 43290 10350 43320
rect 10020 43230 10350 43290
rect 9780 43050 9840 43230
rect 10290 43110 10350 43230
rect 9600 42990 9840 43050
rect 9330 42570 9390 42690
rect 9330 42510 9420 42570
rect 9360 42480 9420 42510
rect 9510 42480 9570 42930
rect 10020 42720 10080 42990
rect 9870 42660 10080 42720
rect 9870 42480 9930 42660
rect 10290 42570 10350 42990
rect 11010 42690 11070 43620
rect 10980 42570 11070 42690
rect 11250 43530 11310 43620
rect 11250 43410 11340 43530
rect 10020 42510 10350 42570
rect 11010 42510 11160 42570
rect 10020 42480 10080 42510
rect 10290 42480 10350 42510
rect 11100 42480 11160 42510
rect 11250 42480 11310 43410
rect 12450 42690 12510 43620
rect 12420 42570 12510 42690
rect 12690 43530 12750 43620
rect 12690 43410 12780 43530
rect 12450 42510 12600 42570
rect 12540 42480 12600 42510
rect 12690 42480 12750 43410
rect 21330 43530 21390 43620
rect 21300 43410 21390 43530
rect 13890 43170 13950 43320
rect 13800 42690 13860 43110
rect 14130 42930 14190 43320
rect 14100 42810 14190 42930
rect 13800 42630 13950 42690
rect 13890 42480 13950 42630
rect 14130 42570 14190 42810
rect 14040 42510 14190 42570
rect 14040 42480 14100 42510
rect 7980 41880 8040 42150
rect 14370 42210 14430 43320
rect 15570 43230 15630 43320
rect 15720 43290 15780 43320
rect 15720 43230 15870 43290
rect 15540 43110 15630 43230
rect 14280 41880 14340 42150
rect 15570 41880 15630 43110
rect 15810 42390 15870 43230
rect 17250 43170 17310 43320
rect 17160 42690 17220 43110
rect 17490 42930 17550 43320
rect 17460 42810 17550 42930
rect 17160 42630 17310 42690
rect 17250 42480 17310 42630
rect 17490 42570 17550 42810
rect 17400 42510 17550 42570
rect 17400 42480 17460 42510
rect 15810 42270 15900 42390
rect 15810 41880 15870 42270
rect 17730 42210 17790 43320
rect 19410 43290 19470 43320
rect 19680 43290 19740 43320
rect 19410 43230 19740 43290
rect 19830 43290 19890 43320
rect 20190 43290 20250 43320
rect 19830 43230 19980 43290
rect 19410 43110 19470 43230
rect 19920 43050 19980 43230
rect 20220 43230 20250 43290
rect 20340 43290 20400 43320
rect 20340 43230 20460 43290
rect 19920 42990 20130 43050
rect 19410 42570 19470 42990
rect 19740 42900 19800 42990
rect 19740 42840 19890 42900
rect 19410 42510 19740 42570
rect 19410 42480 19470 42510
rect 19680 42480 19740 42510
rect 19830 42480 19890 42840
rect 20070 42690 20130 42990
rect 20400 42870 20460 43230
rect 20610 43110 20670 43320
rect 20190 42480 20250 42690
rect 20400 42570 20460 42750
rect 20640 42600 20700 42990
rect 20340 42510 20460 42570
rect 20610 42540 20700 42600
rect 20340 42480 20400 42510
rect 20610 42480 20670 42540
rect 17640 41880 17700 42150
rect 21330 41880 21390 43410
rect 34770 43530 34830 43620
rect 34740 43410 34830 43530
rect 22770 43110 22830 43320
rect 23040 43290 23100 43320
rect 22980 43230 23100 43290
rect 23190 43290 23250 43320
rect 23550 43290 23610 43320
rect 22770 42480 22830 42990
rect 22980 42810 23040 43230
rect 23190 43170 23220 43290
rect 23460 43230 23610 43290
rect 23700 43290 23760 43320
rect 23970 43290 24030 43320
rect 23700 43230 24030 43290
rect 23460 43050 23520 43230
rect 23970 43110 24030 43230
rect 23280 42990 23520 43050
rect 23010 42570 23070 42690
rect 23010 42510 23100 42570
rect 23040 42480 23100 42510
rect 23190 42480 23250 42930
rect 23700 42720 23760 42990
rect 23550 42660 23760 42720
rect 23550 42480 23610 42660
rect 23970 42570 24030 42990
rect 23700 42510 24030 42570
rect 23700 42480 23760 42510
rect 23970 42480 24030 42510
rect 25170 42210 25230 43320
rect 25410 42930 25470 43320
rect 25650 43170 25710 43320
rect 26850 43230 26910 43320
rect 27000 43290 27060 43320
rect 27000 43230 27150 43290
rect 26820 43110 26910 43230
rect 25410 42810 25500 42930
rect 25410 42570 25470 42810
rect 25740 42690 25800 43110
rect 25650 42630 25800 42690
rect 25410 42510 25560 42570
rect 25500 42480 25560 42510
rect 25650 42480 25710 42630
rect 25260 41880 25320 42150
rect 26850 41880 26910 43110
rect 27090 42390 27150 43230
rect 28050 43170 28110 43320
rect 27960 42690 28020 43110
rect 28290 42930 28350 43320
rect 28260 42810 28350 42930
rect 27960 42630 28110 42690
rect 28050 42480 28110 42630
rect 28290 42570 28350 42810
rect 28200 42510 28350 42570
rect 28200 42480 28260 42510
rect 27090 42270 27180 42390
rect 27090 41880 27150 42270
rect 28530 42210 28590 43320
rect 29250 43230 29310 43320
rect 29400 43290 29460 43320
rect 29400 43230 29550 43290
rect 29220 43110 29310 43230
rect 28440 41880 28500 42150
rect 29250 41880 29310 43110
rect 29490 42390 29550 43230
rect 30450 43170 30510 43320
rect 30360 42690 30420 43110
rect 30690 42930 30750 43320
rect 30660 42810 30750 42930
rect 30360 42630 30510 42690
rect 30450 42480 30510 42630
rect 30690 42570 30750 42810
rect 30600 42510 30750 42570
rect 30600 42480 30660 42510
rect 29490 42270 29580 42390
rect 29490 41880 29550 42270
rect 30930 42210 30990 43320
rect 31890 43170 31950 43320
rect 31800 42690 31860 43110
rect 32130 42930 32190 43320
rect 32100 42810 32190 42930
rect 31800 42630 31950 42690
rect 31890 42480 31950 42630
rect 32130 42570 32190 42810
rect 32040 42510 32190 42570
rect 32040 42480 32100 42510
rect 30840 41880 30900 42150
rect 32370 42210 32430 43320
rect 33420 43290 33480 43320
rect 33330 43230 33480 43290
rect 33570 43230 33630 43320
rect 33330 42390 33390 43230
rect 33300 42270 33390 42390
rect 32280 41880 32340 42150
rect 33330 41880 33390 42270
rect 33570 43110 33660 43230
rect 33570 41880 33630 43110
rect 34770 42480 34830 43410
rect 35010 42690 35070 43620
rect 41970 43530 42030 43620
rect 41940 43410 42030 43530
rect 35970 43110 36030 43320
rect 36240 43290 36300 43320
rect 36180 43230 36300 43290
rect 36390 43290 36450 43320
rect 36750 43290 36810 43320
rect 35010 42570 35100 42690
rect 34920 42510 35070 42570
rect 34920 42480 34980 42510
rect 35970 42480 36030 42990
rect 36180 42810 36240 43230
rect 36390 43170 36420 43290
rect 36660 43230 36810 43290
rect 36900 43290 36960 43320
rect 37170 43290 37230 43320
rect 36900 43230 37230 43290
rect 36660 43050 36720 43230
rect 37170 43110 37230 43230
rect 36480 42990 36720 43050
rect 36210 42570 36270 42690
rect 36210 42510 36300 42570
rect 36240 42480 36300 42510
rect 36390 42480 36450 42930
rect 36900 42720 36960 42990
rect 36750 42660 36960 42720
rect 36750 42480 36810 42660
rect 37170 42570 37230 42990
rect 36900 42510 37230 42570
rect 36900 42480 36960 42510
rect 37170 42480 37230 42510
rect 37890 42210 37950 43320
rect 38130 42930 38190 43320
rect 38370 43170 38430 43320
rect 39570 43290 39630 43320
rect 39840 43290 39900 43320
rect 39570 43230 39900 43290
rect 39990 43290 40050 43320
rect 40350 43290 40410 43320
rect 39990 43230 40140 43290
rect 39570 43110 39630 43230
rect 38130 42810 38220 42930
rect 38130 42570 38190 42810
rect 38460 42690 38520 43110
rect 40080 43050 40140 43230
rect 40380 43170 40410 43290
rect 40500 43290 40560 43320
rect 40500 43230 40620 43290
rect 40080 42990 40320 43050
rect 38370 42630 38520 42690
rect 38130 42510 38280 42570
rect 38220 42480 38280 42510
rect 38370 42480 38430 42630
rect 39570 42570 39630 42990
rect 39840 42720 39900 42990
rect 39840 42660 40050 42720
rect 39570 42510 39900 42570
rect 39570 42480 39630 42510
rect 39840 42480 39900 42510
rect 39990 42480 40050 42660
rect 40350 42480 40410 42930
rect 40560 42810 40620 43230
rect 40770 43110 40830 43320
rect 40530 42570 40590 42690
rect 40500 42510 40590 42570
rect 40500 42480 40560 42510
rect 40770 42480 40830 42990
rect 37980 41880 38040 42150
rect 41970 41880 42030 43410
rect 45330 43530 45390 43620
rect 45330 43410 45420 43530
rect 43170 43170 43230 43320
rect 43080 42690 43140 43110
rect 43410 42930 43470 43320
rect 43380 42810 43470 42930
rect 43080 42630 43230 42690
rect 43170 42480 43230 42630
rect 43410 42570 43470 42810
rect 43320 42510 43470 42570
rect 43320 42480 43380 42510
rect 43650 42210 43710 43320
rect 44370 43170 44430 43320
rect 44280 42690 44340 43110
rect 44610 42930 44670 43320
rect 44580 42810 44670 42930
rect 44280 42630 44430 42690
rect 44370 42480 44430 42630
rect 44610 42570 44670 42810
rect 44520 42510 44670 42570
rect 44520 42480 44580 42510
rect 43560 41880 43620 42150
rect 44850 42210 44910 43320
rect 44760 41880 44820 42150
rect 45330 41880 45390 43410
rect 45810 43110 45870 43320
rect 46080 43290 46140 43320
rect 46020 43230 46140 43290
rect 46230 43290 46290 43320
rect 46590 43290 46650 43320
rect 45810 42480 45870 42990
rect 46020 42810 46080 43230
rect 46230 43170 46260 43290
rect 46500 43230 46650 43290
rect 46740 43290 46800 43320
rect 47010 43290 47070 43320
rect 46740 43230 47070 43290
rect 46500 43050 46560 43230
rect 47010 43110 47070 43230
rect 47490 43110 47550 43320
rect 47760 43290 47820 43320
rect 47700 43230 47820 43290
rect 47910 43290 47970 43320
rect 48270 43290 48330 43320
rect 46320 42990 46560 43050
rect 46050 42570 46110 42690
rect 46050 42510 46140 42570
rect 46080 42480 46140 42510
rect 46230 42480 46290 42930
rect 46740 42720 46800 42990
rect 46590 42660 46800 42720
rect 46590 42480 46650 42660
rect 47010 42570 47070 42990
rect 46740 42510 47070 42570
rect 46740 42480 46800 42510
rect 47010 42480 47070 42510
rect 47490 42480 47550 42990
rect 47700 42810 47760 43230
rect 47910 43170 47940 43290
rect 48180 43230 48330 43290
rect 48420 43290 48480 43320
rect 48690 43290 48750 43320
rect 48420 43230 48750 43290
rect 48180 43050 48240 43230
rect 48690 43110 48750 43230
rect 48000 42990 48240 43050
rect 47730 42570 47790 42690
rect 47730 42510 47820 42570
rect 47760 42480 47820 42510
rect 47910 42480 47970 42930
rect 48420 42720 48480 42990
rect 48270 42660 48480 42720
rect 48270 42480 48330 42660
rect 48690 42570 48750 42990
rect 48420 42510 48750 42570
rect 48420 42480 48480 42510
rect 48690 42480 48750 42510
rect 5820 41220 5880 41280
rect 6060 41220 6120 41280
rect 6210 41220 6270 41280
rect 6930 41220 6990 41280
rect 7170 41220 7230 41280
rect 7980 41220 8040 41280
rect 8220 41220 8280 41280
rect 8370 41220 8430 41280
rect 9090 41220 9150 41280
rect 9360 41220 9420 41280
rect 9510 41220 9570 41280
rect 9870 41220 9930 41280
rect 10020 41220 10080 41280
rect 10290 41220 10350 41280
rect 11100 41220 11160 41280
rect 11250 41220 11310 41280
rect 12540 41220 12600 41280
rect 12690 41220 12750 41280
rect 13890 41220 13950 41280
rect 14040 41220 14100 41280
rect 14280 41220 14340 41280
rect 15570 41220 15630 41280
rect 15810 41220 15870 41280
rect 17250 41220 17310 41280
rect 17400 41220 17460 41280
rect 17640 41220 17700 41280
rect 19410 41220 19470 41280
rect 19680 41220 19740 41280
rect 19830 41220 19890 41280
rect 20190 41220 20250 41280
rect 20340 41220 20400 41280
rect 20610 41220 20670 41280
rect 21330 41220 21390 41280
rect 22770 41220 22830 41280
rect 23040 41220 23100 41280
rect 23190 41220 23250 41280
rect 23550 41220 23610 41280
rect 23700 41220 23760 41280
rect 23970 41220 24030 41280
rect 25260 41220 25320 41280
rect 25500 41220 25560 41280
rect 25650 41220 25710 41280
rect 26850 41220 26910 41280
rect 27090 41220 27150 41280
rect 28050 41220 28110 41280
rect 28200 41220 28260 41280
rect 28440 41220 28500 41280
rect 29250 41220 29310 41280
rect 29490 41220 29550 41280
rect 30450 41220 30510 41280
rect 30600 41220 30660 41280
rect 30840 41220 30900 41280
rect 31890 41220 31950 41280
rect 32040 41220 32100 41280
rect 32280 41220 32340 41280
rect 33330 41220 33390 41280
rect 33570 41220 33630 41280
rect 34770 41220 34830 41280
rect 34920 41220 34980 41280
rect 35970 41220 36030 41280
rect 36240 41220 36300 41280
rect 36390 41220 36450 41280
rect 36750 41220 36810 41280
rect 36900 41220 36960 41280
rect 37170 41220 37230 41280
rect 37980 41220 38040 41280
rect 38220 41220 38280 41280
rect 38370 41220 38430 41280
rect 39570 41220 39630 41280
rect 39840 41220 39900 41280
rect 39990 41220 40050 41280
rect 40350 41220 40410 41280
rect 40500 41220 40560 41280
rect 40770 41220 40830 41280
rect 41970 41220 42030 41280
rect 43170 41220 43230 41280
rect 43320 41220 43380 41280
rect 43560 41220 43620 41280
rect 44370 41220 44430 41280
rect 44520 41220 44580 41280
rect 44760 41220 44820 41280
rect 45330 41220 45390 41280
rect 45810 41220 45870 41280
rect 46080 41220 46140 41280
rect 46230 41220 46290 41280
rect 46590 41220 46650 41280
rect 46740 41220 46800 41280
rect 47010 41220 47070 41280
rect 47490 41220 47550 41280
rect 47760 41220 47820 41280
rect 47910 41220 47970 41280
rect 48270 41220 48330 41280
rect 48420 41220 48480 41280
rect 48690 41220 48750 41280
rect 5970 40920 6030 40980
rect 6210 40920 6270 40980
rect 6450 40920 6510 40980
rect 8370 40920 8430 40980
rect 8610 40920 8670 40980
rect 9810 40920 9870 40980
rect 10050 40920 10110 40980
rect 10770 40920 10830 40980
rect 11010 40920 11070 40980
rect 11250 40920 11310 40980
rect 11730 40920 11790 40980
rect 12000 40920 12060 40980
rect 12150 40920 12210 40980
rect 12510 40920 12570 40980
rect 12660 40920 12720 40980
rect 12930 40920 12990 40980
rect 13650 40920 13710 40980
rect 13890 40920 13950 40980
rect 14610 40920 14670 40980
rect 14850 40920 14910 40980
rect 15090 40920 15150 40980
rect 15810 40920 15870 40980
rect 16530 40920 16590 40980
rect 16680 40920 16740 40980
rect 16920 40920 16980 40980
rect 17820 40920 17880 40980
rect 18060 40920 18120 40980
rect 18210 40920 18270 40980
rect 18690 40920 18750 40980
rect 19410 40920 19470 40980
rect 19560 40920 19620 40980
rect 19800 40920 19860 40980
rect 21090 40920 21150 40980
rect 21330 40920 21390 40980
rect 22050 40920 22110 40980
rect 22320 40920 22380 40980
rect 22470 40920 22530 40980
rect 22830 40920 22890 40980
rect 22980 40920 23040 40980
rect 23250 40920 23310 40980
rect 23970 40920 24030 40980
rect 24120 40920 24180 40980
rect 24930 40920 24990 40980
rect 25080 40920 25140 40980
rect 25320 40920 25380 40980
rect 26370 40920 26430 40980
rect 26610 40920 26670 40980
rect 26850 40920 26910 40980
rect 27090 40920 27150 40980
rect 28050 40920 28110 40980
rect 30690 40920 30750 40980
rect 30930 40920 30990 40980
rect 32130 40920 32190 40980
rect 32370 40920 32430 40980
rect 33570 40920 33630 40980
rect 33840 40920 33900 40980
rect 33990 40920 34050 40980
rect 34350 40920 34410 40980
rect 34500 40920 34560 40980
rect 34770 40920 34830 40980
rect 36210 40920 36270 40980
rect 36360 40920 36420 40980
rect 36600 40920 36660 40980
rect 37890 40920 37950 40980
rect 38130 40920 38190 40980
rect 39090 40920 39150 40980
rect 39240 40920 39300 40980
rect 39480 40920 39540 40980
rect 40530 40920 40590 40980
rect 40770 40920 40830 40980
rect 41970 40920 42030 40980
rect 43170 40920 43230 40980
rect 43320 40920 43380 40980
rect 43560 40920 43620 40980
rect 44850 40920 44910 40980
rect 46140 40920 46200 40980
rect 46380 40920 46440 40980
rect 46530 40920 46590 40980
rect 47730 40920 47790 40980
rect 47880 40920 47940 40980
rect 48120 40920 48180 40980
rect 49410 40920 49470 40980
rect 49650 40920 49710 40980
rect 8370 39930 8430 40320
rect 8340 39810 8430 39930
rect 5970 39570 6030 39720
rect 5880 38970 5940 39510
rect 6210 39330 6270 39720
rect 6180 39210 6270 39330
rect 5880 38910 6120 38970
rect 6060 38880 6120 38910
rect 6210 38880 6270 39210
rect 6450 38580 6510 39720
rect 8370 38970 8430 39810
rect 8610 39090 8670 40320
rect 9810 39090 9870 40320
rect 8610 38970 8700 39090
rect 9780 38970 9870 39090
rect 10050 39930 10110 40320
rect 10050 39810 10140 39930
rect 10050 38970 10110 39810
rect 8370 38910 8520 38970
rect 8460 38880 8520 38910
rect 8610 38880 8670 38970
rect 9810 38880 9870 38970
rect 9960 38910 10110 38970
rect 9960 38880 10020 38910
rect 10770 38580 10830 39720
rect 11010 39330 11070 39720
rect 11250 39570 11310 39720
rect 11730 39660 11790 39720
rect 12000 39690 12060 39720
rect 11700 39600 11790 39660
rect 11940 39630 12060 39690
rect 11010 39210 11100 39330
rect 11010 38880 11070 39210
rect 11340 38970 11400 39510
rect 11700 39210 11760 39600
rect 11940 39450 12000 39630
rect 12150 39510 12210 39720
rect 11160 38910 11400 38970
rect 11160 38880 11220 38910
rect 11730 38880 11790 39090
rect 11940 38970 12000 39330
rect 12270 39210 12330 39510
rect 12510 39360 12570 39720
rect 12660 39690 12720 39720
rect 12930 39690 12990 39720
rect 12660 39630 12990 39690
rect 12510 39300 12660 39360
rect 12600 39210 12660 39300
rect 12930 39210 12990 39630
rect 12270 39150 12480 39210
rect 11940 38910 12060 38970
rect 12000 38880 12060 38910
rect 12150 38910 12180 38970
rect 12420 38970 12480 39150
rect 13650 39090 13710 40320
rect 12930 38970 12990 39090
rect 13620 38970 13710 39090
rect 13890 39930 13950 40320
rect 13890 39810 13980 39930
rect 13890 38970 13950 39810
rect 14610 39090 14670 40320
rect 14850 39690 14910 40320
rect 14850 39270 14910 39570
rect 15090 39330 15150 40320
rect 14850 39210 15000 39270
rect 14610 39000 14640 39090
rect 12420 38910 12570 38970
rect 12150 38880 12210 38910
rect 12510 38880 12570 38910
rect 12660 38910 12990 38970
rect 12660 38880 12720 38910
rect 12930 38880 12990 38910
rect 13650 38880 13710 38970
rect 13800 38910 13950 38970
rect 13800 38880 13860 38910
rect 14700 38580 14760 38970
rect 14940 38880 15000 39210
rect 15090 39210 15180 39330
rect 15090 38880 15150 39210
rect 15810 38790 15870 40320
rect 16920 40050 16980 40320
rect 17820 40050 17880 40320
rect 16530 39570 16590 39720
rect 16680 39690 16740 39720
rect 16680 39630 16830 39690
rect 16440 39510 16590 39570
rect 16440 39090 16500 39510
rect 16770 39390 16830 39630
rect 16740 39270 16830 39390
rect 16530 38880 16590 39030
rect 16770 38880 16830 39270
rect 17010 38880 17070 39990
rect 17730 38880 17790 39990
rect 18060 39690 18120 39720
rect 17970 39630 18120 39690
rect 17970 39390 18030 39630
rect 18210 39570 18270 39720
rect 18210 39510 18360 39570
rect 17970 39270 18060 39390
rect 17970 38880 18030 39270
rect 18300 39090 18360 39510
rect 18210 38880 18270 39030
rect 15780 38670 15870 38790
rect 15810 38580 15870 38670
rect 18690 38790 18750 40320
rect 19800 40050 19860 40320
rect 19410 39570 19470 39720
rect 19560 39690 19620 39720
rect 19560 39630 19710 39690
rect 19320 39510 19470 39570
rect 19320 39090 19380 39510
rect 19650 39390 19710 39630
rect 19620 39270 19710 39390
rect 19410 38880 19470 39030
rect 19650 38880 19710 39270
rect 19890 38880 19950 39990
rect 21090 39930 21150 40320
rect 21060 39810 21150 39930
rect 21090 38970 21150 39810
rect 21330 39090 21390 40320
rect 25320 40050 25380 40320
rect 22050 39210 22110 39720
rect 22320 39690 22380 39720
rect 22290 39630 22380 39690
rect 22290 39510 22350 39630
rect 21330 38970 21420 39090
rect 21090 38910 21240 38970
rect 21180 38880 21240 38910
rect 21330 38880 21390 38970
rect 22050 38880 22110 39090
rect 22260 38970 22320 39390
rect 22470 39270 22530 39720
rect 22830 39540 22890 39720
rect 22980 39690 23040 39720
rect 23250 39690 23310 39720
rect 22980 39630 23310 39690
rect 22830 39480 23040 39540
rect 22980 39210 23040 39480
rect 23250 39210 23310 39630
rect 22560 39150 22800 39210
rect 22260 38910 22380 38970
rect 22320 38880 22380 38910
rect 22470 38910 22500 39030
rect 22740 38970 22800 39150
rect 23250 38970 23310 39090
rect 22740 38910 22890 38970
rect 22470 38880 22530 38910
rect 22830 38880 22890 38910
rect 22980 38910 23310 38970
rect 22980 38880 23040 38910
rect 23250 38880 23310 38910
rect 18690 38670 18780 38790
rect 18690 38580 18750 38670
rect 23970 38790 24030 39720
rect 24120 39690 24180 39720
rect 24120 39630 24270 39690
rect 23940 38670 24030 38790
rect 23970 38580 24030 38670
rect 24210 39510 24300 39630
rect 24930 39570 24990 39720
rect 25080 39690 25140 39720
rect 25080 39630 25230 39690
rect 24840 39510 24990 39570
rect 24210 38580 24270 39510
rect 24840 39090 24900 39510
rect 25170 39390 25230 39630
rect 25140 39270 25230 39390
rect 24930 38880 24990 39030
rect 25170 38880 25230 39270
rect 25410 38880 25470 39990
rect 26370 39570 26430 39720
rect 26610 39690 26670 39720
rect 26580 39630 26670 39690
rect 26280 38970 26340 39510
rect 26280 38910 26490 38970
rect 26430 38880 26490 38910
rect 26580 38880 26640 39630
rect 26850 39300 26910 39720
rect 27090 39690 27150 39720
rect 27090 39630 27210 39690
rect 27150 39510 27180 39630
rect 26880 39270 26910 39300
rect 26880 38970 26940 39270
rect 27150 39030 27210 39510
rect 27090 38970 27210 39030
rect 26880 38910 27000 38970
rect 26940 38880 27000 38910
rect 27090 38880 27150 38970
rect 28050 38790 28110 40320
rect 30690 39930 30750 40320
rect 30660 39810 30750 39930
rect 30690 38970 30750 39810
rect 30930 39090 30990 40320
rect 32130 39930 32190 40320
rect 32100 39810 32190 39930
rect 30930 38970 31020 39090
rect 32130 38970 32190 39810
rect 32370 39090 32430 40320
rect 36600 40050 36660 40320
rect 33570 39210 33630 39720
rect 33840 39690 33900 39720
rect 33810 39630 33900 39690
rect 33810 39510 33870 39630
rect 32370 38970 32460 39090
rect 30690 38910 30840 38970
rect 30780 38880 30840 38910
rect 30930 38880 30990 38970
rect 32130 38910 32280 38970
rect 32220 38880 32280 38910
rect 32370 38880 32430 38970
rect 33570 38880 33630 39090
rect 33780 38970 33840 39390
rect 33990 39270 34050 39720
rect 34350 39540 34410 39720
rect 34500 39690 34560 39720
rect 34770 39690 34830 39720
rect 34500 39630 34830 39690
rect 34350 39480 34560 39540
rect 34500 39210 34560 39480
rect 34770 39210 34830 39630
rect 36210 39570 36270 39720
rect 36360 39690 36420 39720
rect 36360 39630 36510 39690
rect 36120 39510 36270 39570
rect 34080 39150 34320 39210
rect 33780 38910 33900 38970
rect 33840 38880 33900 38910
rect 33990 38910 34020 39030
rect 34260 38970 34320 39150
rect 36120 39090 36180 39510
rect 36450 39390 36510 39630
rect 36420 39270 36510 39390
rect 34770 38970 34830 39090
rect 34260 38910 34410 38970
rect 33990 38880 34050 38910
rect 34350 38880 34410 38910
rect 34500 38910 34830 38970
rect 34500 38880 34560 38910
rect 34770 38880 34830 38910
rect 36210 38880 36270 39030
rect 36450 38880 36510 39270
rect 36690 38880 36750 39990
rect 37890 39930 37950 40320
rect 37860 39810 37950 39930
rect 37890 38970 37950 39810
rect 38130 39090 38190 40320
rect 39480 40050 39540 40320
rect 39090 39570 39150 39720
rect 39240 39690 39300 39720
rect 39240 39630 39390 39690
rect 39000 39510 39150 39570
rect 39000 39090 39060 39510
rect 39330 39390 39390 39630
rect 39300 39270 39390 39390
rect 38130 38970 38220 39090
rect 37890 38910 38040 38970
rect 37980 38880 38040 38910
rect 38130 38880 38190 38970
rect 39090 38880 39150 39030
rect 39330 38880 39390 39270
rect 39570 38880 39630 39990
rect 40530 39090 40590 40320
rect 40500 38970 40590 39090
rect 40770 39930 40830 40320
rect 40770 39810 40860 39930
rect 40770 38970 40830 39810
rect 40530 38880 40590 38970
rect 40680 38910 40830 38970
rect 40680 38880 40740 38910
rect 28050 38670 28140 38790
rect 28050 38580 28110 38670
rect 41970 38790 42030 40320
rect 43560 40050 43620 40320
rect 43170 39570 43230 39720
rect 43320 39690 43380 39720
rect 43320 39630 43470 39690
rect 43080 39510 43230 39570
rect 43080 39090 43140 39510
rect 43410 39390 43470 39630
rect 43380 39270 43470 39390
rect 43170 38880 43230 39030
rect 43410 38880 43470 39270
rect 43650 38880 43710 39990
rect 41940 38670 42030 38790
rect 41970 38580 42030 38670
rect 44850 38790 44910 40320
rect 46140 40050 46200 40320
rect 46050 38880 46110 39990
rect 48120 40050 48180 40320
rect 46380 39690 46440 39720
rect 46290 39630 46440 39690
rect 46290 39390 46350 39630
rect 46530 39570 46590 39720
rect 47730 39570 47790 39720
rect 47880 39690 47940 39720
rect 47880 39630 48030 39690
rect 46530 39510 46680 39570
rect 46290 39270 46380 39390
rect 46290 38880 46350 39270
rect 46620 39090 46680 39510
rect 47640 39510 47790 39570
rect 47640 39090 47700 39510
rect 47970 39390 48030 39630
rect 47940 39270 48030 39390
rect 46530 38880 46590 39030
rect 47730 38880 47790 39030
rect 47970 38880 48030 39270
rect 48210 38880 48270 39990
rect 49410 39930 49470 40320
rect 49380 39810 49470 39930
rect 49410 38970 49470 39810
rect 49650 39090 49710 40320
rect 49650 38970 49740 39090
rect 49410 38910 49560 38970
rect 49500 38880 49560 38910
rect 49650 38880 49710 38970
rect 44820 38670 44910 38790
rect 44850 38580 44910 38670
rect 6060 38220 6120 38280
rect 6210 38220 6270 38280
rect 6450 38220 6510 38280
rect 8460 38220 8520 38280
rect 8610 38220 8670 38280
rect 9810 38220 9870 38280
rect 9960 38220 10020 38280
rect 10770 38220 10830 38280
rect 11010 38220 11070 38280
rect 11160 38220 11220 38280
rect 11730 38220 11790 38280
rect 12000 38220 12060 38280
rect 12150 38220 12210 38280
rect 12510 38220 12570 38280
rect 12660 38220 12720 38280
rect 12930 38220 12990 38280
rect 13650 38220 13710 38280
rect 13800 38220 13860 38280
rect 14700 38220 14760 38280
rect 14940 38220 15000 38280
rect 15090 38220 15150 38280
rect 15810 38220 15870 38280
rect 16530 38220 16590 38280
rect 16770 38220 16830 38280
rect 17010 38220 17070 38280
rect 17730 38220 17790 38280
rect 17970 38220 18030 38280
rect 18210 38220 18270 38280
rect 18690 38220 18750 38280
rect 19410 38220 19470 38280
rect 19650 38220 19710 38280
rect 19890 38220 19950 38280
rect 21180 38220 21240 38280
rect 21330 38220 21390 38280
rect 22050 38220 22110 38280
rect 22320 38220 22380 38280
rect 22470 38220 22530 38280
rect 22830 38220 22890 38280
rect 22980 38220 23040 38280
rect 23250 38220 23310 38280
rect 23970 38220 24030 38280
rect 24210 38220 24270 38280
rect 24930 38220 24990 38280
rect 25170 38220 25230 38280
rect 25410 38220 25470 38280
rect 26430 38220 26490 38280
rect 26580 38220 26640 38280
rect 26940 38220 27000 38280
rect 27090 38220 27150 38280
rect 28050 38220 28110 38280
rect 30780 38220 30840 38280
rect 30930 38220 30990 38280
rect 32220 38220 32280 38280
rect 32370 38220 32430 38280
rect 33570 38220 33630 38280
rect 33840 38220 33900 38280
rect 33990 38220 34050 38280
rect 34350 38220 34410 38280
rect 34500 38220 34560 38280
rect 34770 38220 34830 38280
rect 36210 38220 36270 38280
rect 36450 38220 36510 38280
rect 36690 38220 36750 38280
rect 37980 38220 38040 38280
rect 38130 38220 38190 38280
rect 39090 38220 39150 38280
rect 39330 38220 39390 38280
rect 39570 38220 39630 38280
rect 40530 38220 40590 38280
rect 40680 38220 40740 38280
rect 41970 38220 42030 38280
rect 43170 38220 43230 38280
rect 43410 38220 43470 38280
rect 43650 38220 43710 38280
rect 44850 38220 44910 38280
rect 46050 38220 46110 38280
rect 46290 38220 46350 38280
rect 46530 38220 46590 38280
rect 47730 38220 47790 38280
rect 47970 38220 48030 38280
rect 48210 38220 48270 38280
rect 49500 38220 49560 38280
rect 49650 38220 49710 38280
rect 5820 37920 5880 37980
rect 5970 37920 6030 37980
rect 7170 37920 7230 37980
rect 8370 37920 8430 37980
rect 8610 37920 8670 37980
rect 8850 37920 8910 37980
rect 11010 37920 11070 37980
rect 11160 37920 11220 37980
rect 12210 37920 12270 37980
rect 12450 37920 12510 37980
rect 12690 37920 12750 37980
rect 15090 37920 15150 37980
rect 15330 37920 15390 37980
rect 15570 37920 15630 37980
rect 16860 37920 16920 37980
rect 17100 37920 17160 37980
rect 17250 37920 17310 37980
rect 18210 37920 18270 37980
rect 18360 37920 18420 37980
rect 19650 37920 19710 37980
rect 19800 37920 19860 37980
rect 21090 37920 21150 37980
rect 21240 37920 21300 37980
rect 22530 37920 22590 37980
rect 22680 37920 22740 37980
rect 23970 37920 24030 37980
rect 25260 37920 25320 37980
rect 25410 37920 25470 37980
rect 26610 37920 26670 37980
rect 26850 37920 26910 37980
rect 27090 37920 27150 37980
rect 28050 37920 28110 37980
rect 28200 37920 28260 37980
rect 29250 37920 29310 37980
rect 29400 37920 29460 37980
rect 30210 37920 30270 37980
rect 30450 37920 30510 37980
rect 30690 37920 30750 37980
rect 31410 37920 31470 37980
rect 32130 37920 32190 37980
rect 32370 37920 32430 37980
rect 32610 37920 32670 37980
rect 33420 37920 33480 37980
rect 33570 37920 33630 37980
rect 34770 37920 34830 37980
rect 34920 37920 34980 37980
rect 35730 37920 35790 37980
rect 36000 37920 36060 37980
rect 36150 37920 36210 37980
rect 36510 37920 36570 37980
rect 36660 37920 36720 37980
rect 36930 37920 36990 37980
rect 39090 37920 39150 37980
rect 40050 37920 40110 37980
rect 40200 37920 40260 37980
rect 40560 37920 40620 37980
rect 40710 37920 40770 37980
rect 41730 37920 41790 37980
rect 42450 37920 42510 37980
rect 42690 37920 42750 37980
rect 42930 37920 42990 37980
rect 43650 37920 43710 37980
rect 44610 37920 44670 37980
rect 44850 37920 44910 37980
rect 45090 37920 45150 37980
rect 46290 37920 46350 37980
rect 46440 37920 46500 37980
rect 47730 37920 47790 37980
rect 47970 37920 48030 37980
rect 48210 37920 48270 37980
rect 49500 37920 49560 37980
rect 49650 37920 49710 37980
rect 7170 37530 7230 37620
rect 7170 37410 7260 37530
rect 5820 37290 5880 37320
rect 5730 37230 5880 37290
rect 5970 37230 6030 37320
rect 5730 36390 5790 37230
rect 5700 36270 5790 36390
rect 5730 35880 5790 36270
rect 5970 37110 6060 37230
rect 5970 35880 6030 37110
rect 7170 35880 7230 37410
rect 8370 36210 8430 37320
rect 8610 36930 8670 37320
rect 8850 37170 8910 37320
rect 11010 37230 11070 37320
rect 11160 37290 11220 37320
rect 11160 37230 11310 37290
rect 10980 37110 11070 37230
rect 8610 36810 8700 36930
rect 8610 36570 8670 36810
rect 8940 36690 9000 37110
rect 8850 36630 9000 36690
rect 8610 36510 8760 36570
rect 8700 36480 8760 36510
rect 8850 36480 8910 36630
rect 8460 35880 8520 36150
rect 11010 35880 11070 37110
rect 11250 36390 11310 37230
rect 11250 36270 11340 36390
rect 11250 35880 11310 36270
rect 12210 36210 12270 37320
rect 12450 36930 12510 37320
rect 12690 37170 12750 37320
rect 12450 36810 12540 36930
rect 12450 36570 12510 36810
rect 12780 36690 12840 37110
rect 12690 36630 12840 36690
rect 12450 36510 12600 36570
rect 12540 36480 12600 36510
rect 12690 36480 12750 36630
rect 12300 35880 12360 36150
rect 15090 36210 15150 37320
rect 15330 36930 15390 37320
rect 15570 37170 15630 37320
rect 16860 37230 16920 37620
rect 23970 37530 24030 37620
rect 23940 37410 24030 37530
rect 16770 37110 16800 37200
rect 15330 36810 15420 36930
rect 15330 36570 15390 36810
rect 15660 36690 15720 37110
rect 15570 36630 15720 36690
rect 15330 36510 15480 36570
rect 15420 36480 15480 36510
rect 15570 36480 15630 36630
rect 15180 35880 15240 36150
rect 16770 35880 16830 37110
rect 17100 36990 17160 37320
rect 17010 36930 17160 36990
rect 17250 36990 17310 37320
rect 18210 37230 18270 37320
rect 18360 37290 18420 37320
rect 18360 37230 18510 37290
rect 19650 37230 19710 37320
rect 19800 37290 19860 37320
rect 19800 37230 19950 37290
rect 21090 37230 21150 37320
rect 21240 37290 21300 37320
rect 21240 37230 21390 37290
rect 22530 37230 22590 37320
rect 22680 37290 22740 37320
rect 22680 37230 22830 37290
rect 18180 37110 18270 37230
rect 17010 36630 17070 36930
rect 17250 36870 17340 36990
rect 17010 35880 17070 36510
rect 17250 35880 17310 36870
rect 18210 35880 18270 37110
rect 18450 36390 18510 37230
rect 19620 37110 19710 37230
rect 18450 36270 18540 36390
rect 18450 35880 18510 36270
rect 19650 35880 19710 37110
rect 19890 36390 19950 37230
rect 21060 37110 21150 37230
rect 19890 36270 19980 36390
rect 19890 35880 19950 36270
rect 21090 35880 21150 37110
rect 21330 36390 21390 37230
rect 22500 37110 22590 37230
rect 21330 36270 21420 36390
rect 21330 35880 21390 36270
rect 22530 35880 22590 37110
rect 22770 36390 22830 37230
rect 22770 36270 22860 36390
rect 22770 35880 22830 36270
rect 23970 35880 24030 37410
rect 31410 37530 31470 37620
rect 31380 37410 31470 37530
rect 25260 37290 25320 37320
rect 25170 37230 25320 37290
rect 25410 37230 25470 37320
rect 25170 36390 25230 37230
rect 25140 36270 25230 36390
rect 25170 35880 25230 36270
rect 25410 37110 25500 37230
rect 26610 37170 26670 37320
rect 25410 35880 25470 37110
rect 26520 36690 26580 37110
rect 26850 36930 26910 37320
rect 26820 36810 26910 36930
rect 26520 36630 26670 36690
rect 26610 36480 26670 36630
rect 26850 36570 26910 36810
rect 26760 36510 26910 36570
rect 26760 36480 26820 36510
rect 27090 36210 27150 37320
rect 28050 37230 28110 37320
rect 28200 37290 28260 37320
rect 28200 37230 28350 37290
rect 29250 37230 29310 37320
rect 29400 37290 29460 37320
rect 29400 37230 29550 37290
rect 28020 37110 28110 37230
rect 27000 35880 27060 36150
rect 28050 35880 28110 37110
rect 28290 36390 28350 37230
rect 29220 37110 29310 37230
rect 28290 36270 28380 36390
rect 28290 35880 28350 36270
rect 29250 35880 29310 37110
rect 29490 36390 29550 37230
rect 30210 37170 30270 37320
rect 30120 36690 30180 37110
rect 30450 36930 30510 37320
rect 30420 36810 30510 36930
rect 30120 36630 30270 36690
rect 30210 36480 30270 36630
rect 30450 36570 30510 36810
rect 30360 36510 30510 36570
rect 30360 36480 30420 36510
rect 29490 36270 29580 36390
rect 29490 35880 29550 36270
rect 30690 36210 30750 37320
rect 30600 35880 30660 36150
rect 31410 35880 31470 37410
rect 39090 37530 39150 37620
rect 39060 37410 39150 37530
rect 32130 36210 32190 37320
rect 32370 36930 32430 37320
rect 32610 37170 32670 37320
rect 33420 37290 33480 37320
rect 33330 37230 33480 37290
rect 33570 37230 33630 37320
rect 34770 37230 34830 37320
rect 34920 37290 34980 37320
rect 35730 37290 35790 37320
rect 36000 37290 36060 37320
rect 34920 37230 35070 37290
rect 32370 36810 32460 36930
rect 32370 36570 32430 36810
rect 32700 36690 32760 37110
rect 32610 36630 32760 36690
rect 32370 36510 32520 36570
rect 32460 36480 32520 36510
rect 32610 36480 32670 36630
rect 32220 35880 32280 36150
rect 33330 36390 33390 37230
rect 33300 36270 33390 36390
rect 33330 35880 33390 36270
rect 33570 37110 33660 37230
rect 34740 37110 34830 37230
rect 33570 35880 33630 37110
rect 34770 35880 34830 37110
rect 35010 36390 35070 37230
rect 35730 37230 36060 37290
rect 36150 37290 36210 37320
rect 36510 37290 36570 37320
rect 36150 37230 36300 37290
rect 35730 37110 35790 37230
rect 36240 37050 36300 37230
rect 36540 37170 36570 37290
rect 36660 37290 36720 37320
rect 36660 37230 36780 37290
rect 36240 36990 36480 37050
rect 35730 36570 35790 36990
rect 36000 36720 36060 36990
rect 36000 36660 36210 36720
rect 35730 36510 36060 36570
rect 35730 36480 35790 36510
rect 36000 36480 36060 36510
rect 36150 36480 36210 36660
rect 36510 36480 36570 36930
rect 36720 36810 36780 37230
rect 36930 37110 36990 37320
rect 36690 36570 36750 36690
rect 36660 36510 36750 36570
rect 36660 36480 36720 36510
rect 36930 36480 36990 36990
rect 35010 36270 35100 36390
rect 35010 35880 35070 36270
rect 39090 35880 39150 37410
rect 41730 37530 41790 37620
rect 41700 37410 41790 37530
rect 40050 37230 40110 37320
rect 40200 37290 40260 37320
rect 40200 37230 40320 37290
rect 39990 37170 40110 37230
rect 39990 36690 40050 37170
rect 40260 36930 40320 37230
rect 40290 36900 40320 36930
rect 40020 36570 40050 36690
rect 39990 36510 40110 36570
rect 40050 36480 40110 36510
rect 40290 36480 40350 36900
rect 40560 36570 40620 37320
rect 40710 37290 40770 37320
rect 40710 37230 40920 37290
rect 40860 36690 40920 37230
rect 40530 36510 40620 36570
rect 40530 36480 40590 36510
rect 40770 36480 40830 36630
rect 41730 35880 41790 37410
rect 43650 37530 43710 37620
rect 43650 37410 43740 37530
rect 42450 36210 42510 37320
rect 42690 36930 42750 37320
rect 42930 37170 42990 37320
rect 42690 36810 42780 36930
rect 42690 36570 42750 36810
rect 43020 36690 43080 37110
rect 42930 36630 43080 36690
rect 42690 36510 42840 36570
rect 42780 36480 42840 36510
rect 42930 36480 42990 36630
rect 42540 35880 42600 36150
rect 43650 35880 43710 37410
rect 44610 37170 44670 37320
rect 44520 36690 44580 37110
rect 44850 36930 44910 37320
rect 44820 36810 44910 36930
rect 44520 36630 44670 36690
rect 44610 36480 44670 36630
rect 44850 36570 44910 36810
rect 44760 36510 44910 36570
rect 44760 36480 44820 36510
rect 45090 36210 45150 37320
rect 46290 37230 46350 37320
rect 46440 37290 46500 37320
rect 46440 37230 46590 37290
rect 46260 37110 46350 37230
rect 45000 35880 45060 36150
rect 46290 35880 46350 37110
rect 46530 36390 46590 37230
rect 47730 37170 47790 37320
rect 47640 36690 47700 37110
rect 47970 36930 48030 37320
rect 47940 36810 48030 36930
rect 47640 36630 47790 36690
rect 47730 36480 47790 36630
rect 47970 36570 48030 36810
rect 47880 36510 48030 36570
rect 47880 36480 47940 36510
rect 46530 36270 46620 36390
rect 46530 35880 46590 36270
rect 48210 36210 48270 37320
rect 49500 37290 49560 37320
rect 49410 37230 49560 37290
rect 49650 37230 49710 37320
rect 49410 36390 49470 37230
rect 49380 36270 49470 36390
rect 48120 35880 48180 36150
rect 49410 35880 49470 36270
rect 49650 37110 49740 37230
rect 49650 35880 49710 37110
rect 5730 35220 5790 35280
rect 5970 35220 6030 35280
rect 7170 35220 7230 35280
rect 8460 35220 8520 35280
rect 8700 35220 8760 35280
rect 8850 35220 8910 35280
rect 11010 35220 11070 35280
rect 11250 35220 11310 35280
rect 12300 35220 12360 35280
rect 12540 35220 12600 35280
rect 12690 35220 12750 35280
rect 15180 35220 15240 35280
rect 15420 35220 15480 35280
rect 15570 35220 15630 35280
rect 16770 35220 16830 35280
rect 17010 35220 17070 35280
rect 17250 35220 17310 35280
rect 18210 35220 18270 35280
rect 18450 35220 18510 35280
rect 19650 35220 19710 35280
rect 19890 35220 19950 35280
rect 21090 35220 21150 35280
rect 21330 35220 21390 35280
rect 22530 35220 22590 35280
rect 22770 35220 22830 35280
rect 23970 35220 24030 35280
rect 25170 35220 25230 35280
rect 25410 35220 25470 35280
rect 26610 35220 26670 35280
rect 26760 35220 26820 35280
rect 27000 35220 27060 35280
rect 28050 35220 28110 35280
rect 28290 35220 28350 35280
rect 29250 35220 29310 35280
rect 29490 35220 29550 35280
rect 30210 35220 30270 35280
rect 30360 35220 30420 35280
rect 30600 35220 30660 35280
rect 31410 35220 31470 35280
rect 32220 35220 32280 35280
rect 32460 35220 32520 35280
rect 32610 35220 32670 35280
rect 33330 35220 33390 35280
rect 33570 35220 33630 35280
rect 34770 35220 34830 35280
rect 35010 35220 35070 35280
rect 35730 35220 35790 35280
rect 36000 35220 36060 35280
rect 36150 35220 36210 35280
rect 36510 35220 36570 35280
rect 36660 35220 36720 35280
rect 36930 35220 36990 35280
rect 39090 35220 39150 35280
rect 40050 35220 40110 35280
rect 40290 35220 40350 35280
rect 40530 35220 40590 35280
rect 40770 35220 40830 35280
rect 41730 35220 41790 35280
rect 42540 35220 42600 35280
rect 42780 35220 42840 35280
rect 42930 35220 42990 35280
rect 43650 35220 43710 35280
rect 44610 35220 44670 35280
rect 44760 35220 44820 35280
rect 45000 35220 45060 35280
rect 46290 35220 46350 35280
rect 46530 35220 46590 35280
rect 47730 35220 47790 35280
rect 47880 35220 47940 35280
rect 48120 35220 48180 35280
rect 49410 35220 49470 35280
rect 49650 35220 49710 35280
rect 6780 34920 6840 34980
rect 7020 34920 7080 34980
rect 7170 34920 7230 34980
rect 7980 34920 8040 34980
rect 8220 34920 8280 34980
rect 8370 34920 8430 34980
rect 9090 34920 9150 34980
rect 9360 34920 9420 34980
rect 9510 34920 9570 34980
rect 9870 34920 9930 34980
rect 10020 34920 10080 34980
rect 10290 34920 10350 34980
rect 11250 34920 11310 34980
rect 11520 34920 11580 34980
rect 11670 34920 11730 34980
rect 12030 34920 12090 34980
rect 12180 34920 12240 34980
rect 12450 34920 12510 34980
rect 13890 34920 13950 34980
rect 15330 34920 15390 34980
rect 15570 34920 15630 34980
rect 16770 34920 16830 34980
rect 16920 34920 16980 34980
rect 17160 34920 17220 34980
rect 19410 34920 19470 34980
rect 19650 34920 19710 34980
rect 20850 34920 20910 34980
rect 21090 34920 21150 34980
rect 21330 34920 21390 34980
rect 23490 34920 23550 34980
rect 23640 34920 23700 34980
rect 23880 34920 23940 34980
rect 24930 34920 24990 34980
rect 25080 34920 25140 34980
rect 25320 34920 25380 34980
rect 26130 34920 26190 34980
rect 26400 34920 26460 34980
rect 26550 34920 26610 34980
rect 26910 34920 26970 34980
rect 27060 34920 27120 34980
rect 27330 34920 27390 34980
rect 30450 34920 30510 34980
rect 31170 34920 31230 34980
rect 31410 34920 31470 34980
rect 32130 34920 32190 34980
rect 32280 34920 32340 34980
rect 32520 34920 32580 34980
rect 33330 34920 33390 34980
rect 33570 34920 33630 34980
rect 34770 34920 34830 34980
rect 35010 34920 35070 34980
rect 36210 34920 36270 34980
rect 36450 34920 36510 34980
rect 37650 34920 37710 34980
rect 37890 34920 37950 34980
rect 39090 34920 39150 34980
rect 39330 34920 39390 34980
rect 40290 34920 40350 34980
rect 40440 34920 40500 34980
rect 40680 34920 40740 34980
rect 41730 34920 41790 34980
rect 41970 34920 42030 34980
rect 43170 34920 43230 34980
rect 43320 34920 43380 34980
rect 43560 34920 43620 34980
rect 44370 34920 44430 34980
rect 44640 34920 44700 34980
rect 44790 34920 44850 34980
rect 45150 34920 45210 34980
rect 45300 34920 45360 34980
rect 45570 34920 45630 34980
rect 46290 34920 46350 34980
rect 46440 34920 46500 34980
rect 46680 34920 46740 34980
rect 47730 34920 47790 34980
rect 47970 34920 48030 34980
rect 49170 34920 49230 34980
rect 49410 34920 49470 34980
rect 6780 34050 6840 34320
rect 6690 32880 6750 33990
rect 7980 34050 8040 34320
rect 7020 33690 7080 33720
rect 6930 33630 7080 33690
rect 6930 33390 6990 33630
rect 7170 33570 7230 33720
rect 7170 33510 7320 33570
rect 6930 33270 7020 33390
rect 6930 32880 6990 33270
rect 7260 33090 7320 33510
rect 7170 32880 7230 33030
rect 7890 32880 7950 33990
rect 8220 33690 8280 33720
rect 8130 33630 8280 33690
rect 8130 33390 8190 33630
rect 8370 33570 8430 33720
rect 9090 33660 9150 33720
rect 9360 33690 9420 33720
rect 9060 33600 9150 33660
rect 9300 33630 9420 33690
rect 8370 33510 8520 33570
rect 8130 33270 8220 33390
rect 8130 32880 8190 33270
rect 8460 33090 8520 33510
rect 9060 33210 9120 33600
rect 9300 33450 9360 33630
rect 9510 33510 9570 33720
rect 8370 32880 8430 33030
rect 9090 32880 9150 33090
rect 9300 32970 9360 33330
rect 9630 33210 9690 33510
rect 9870 33360 9930 33720
rect 10020 33690 10080 33720
rect 10290 33690 10350 33720
rect 10020 33630 10350 33690
rect 11250 33660 11310 33720
rect 11520 33690 11580 33720
rect 9870 33300 10020 33360
rect 9960 33210 10020 33300
rect 10290 33210 10350 33630
rect 11220 33600 11310 33660
rect 11460 33630 11580 33690
rect 11220 33210 11280 33600
rect 11460 33450 11520 33630
rect 11670 33510 11730 33720
rect 9630 33150 9840 33210
rect 9300 32910 9420 32970
rect 9360 32880 9420 32910
rect 9510 32910 9540 32970
rect 9780 32970 9840 33150
rect 10290 32970 10350 33090
rect 9780 32910 9930 32970
rect 9510 32880 9570 32910
rect 9870 32880 9930 32910
rect 10020 32910 10350 32970
rect 10020 32880 10080 32910
rect 10290 32880 10350 32910
rect 11250 32880 11310 33090
rect 11460 32970 11520 33330
rect 11790 33210 11850 33510
rect 12030 33360 12090 33720
rect 12180 33690 12240 33720
rect 12450 33690 12510 33720
rect 12180 33630 12510 33690
rect 12030 33300 12180 33360
rect 12120 33210 12180 33300
rect 12450 33210 12510 33630
rect 11790 33150 12000 33210
rect 11460 32910 11580 32970
rect 11520 32880 11580 32910
rect 11670 32910 11700 32970
rect 11940 32970 12000 33150
rect 12450 32970 12510 33090
rect 11940 32910 12090 32970
rect 11670 32880 11730 32910
rect 12030 32880 12090 32910
rect 12180 32910 12510 32970
rect 12180 32880 12240 32910
rect 12450 32880 12510 32910
rect 13890 32790 13950 34320
rect 15330 33090 15390 34320
rect 15300 32970 15390 33090
rect 15570 33930 15630 34320
rect 15570 33810 15660 33930
rect 15570 32970 15630 33810
rect 17160 34050 17220 34320
rect 16770 33570 16830 33720
rect 16920 33690 16980 33720
rect 16920 33630 17070 33690
rect 16680 33510 16830 33570
rect 16680 33090 16740 33510
rect 17010 33390 17070 33630
rect 16980 33270 17070 33390
rect 15330 32880 15390 32970
rect 15480 32910 15630 32970
rect 15480 32880 15540 32910
rect 16770 32880 16830 33030
rect 17010 32880 17070 33270
rect 17250 32880 17310 33990
rect 19410 33930 19470 34320
rect 19380 33810 19470 33930
rect 19410 32970 19470 33810
rect 19650 33090 19710 34320
rect 20850 33090 20910 34320
rect 21090 33690 21150 34320
rect 21090 33270 21150 33570
rect 21330 33330 21390 34320
rect 23880 34050 23940 34320
rect 23490 33570 23550 33720
rect 23640 33690 23700 33720
rect 23640 33630 23790 33690
rect 23400 33510 23550 33570
rect 21090 33210 21240 33270
rect 19650 32970 19740 33090
rect 20850 33000 20880 33090
rect 19410 32910 19560 32970
rect 19500 32880 19560 32910
rect 19650 32880 19710 32970
rect 13890 32670 13980 32790
rect 13890 32580 13950 32670
rect 20940 32580 21000 32970
rect 21180 32880 21240 33210
rect 21330 33210 21420 33330
rect 21330 32880 21390 33210
rect 23400 33090 23460 33510
rect 23730 33390 23790 33630
rect 23700 33270 23790 33390
rect 23490 32880 23550 33030
rect 23730 32880 23790 33270
rect 23970 32880 24030 33990
rect 25320 34050 25380 34320
rect 24930 33570 24990 33720
rect 25080 33690 25140 33720
rect 25080 33630 25230 33690
rect 24840 33510 24990 33570
rect 24840 33090 24900 33510
rect 25170 33390 25230 33630
rect 25140 33270 25230 33390
rect 24930 32880 24990 33030
rect 25170 32880 25230 33270
rect 25410 32880 25470 33990
rect 26130 33210 26190 33720
rect 26400 33690 26460 33720
rect 26370 33630 26460 33690
rect 26370 33510 26430 33630
rect 26130 32880 26190 33090
rect 26340 32970 26400 33390
rect 26550 33270 26610 33720
rect 26910 33540 26970 33720
rect 27060 33690 27120 33720
rect 27330 33690 27390 33720
rect 27060 33630 27390 33690
rect 26910 33480 27120 33540
rect 27060 33210 27120 33480
rect 27330 33210 27390 33630
rect 26640 33150 26880 33210
rect 26340 32910 26460 32970
rect 26400 32880 26460 32910
rect 26550 32910 26580 33030
rect 26820 32970 26880 33150
rect 27330 32970 27390 33090
rect 26820 32910 26970 32970
rect 26550 32880 26610 32910
rect 26910 32880 26970 32910
rect 27060 32910 27390 32970
rect 27060 32880 27120 32910
rect 27330 32880 27390 32910
rect 30450 32790 30510 34320
rect 31170 33930 31230 34320
rect 31140 33810 31230 33930
rect 31170 32970 31230 33810
rect 31410 33090 31470 34320
rect 32520 34050 32580 34320
rect 32130 33570 32190 33720
rect 32280 33690 32340 33720
rect 32280 33630 32430 33690
rect 32040 33510 32190 33570
rect 32040 33090 32100 33510
rect 32370 33390 32430 33630
rect 32340 33270 32430 33390
rect 31410 32970 31500 33090
rect 31170 32910 31320 32970
rect 31260 32880 31320 32910
rect 31410 32880 31470 32970
rect 32130 32880 32190 33030
rect 32370 32880 32430 33270
rect 32610 32880 32670 33990
rect 33330 33090 33390 34320
rect 33300 32970 33390 33090
rect 33570 33930 33630 34320
rect 33570 33810 33660 33930
rect 33570 32970 33630 33810
rect 34770 33090 34830 34320
rect 34740 32970 34830 33090
rect 35010 33930 35070 34320
rect 35010 33810 35100 33930
rect 35010 32970 35070 33810
rect 36210 33090 36270 34320
rect 36180 32970 36270 33090
rect 36450 33930 36510 34320
rect 37650 33930 37710 34320
rect 36450 33810 36540 33930
rect 37620 33810 37710 33930
rect 36450 32970 36510 33810
rect 33330 32880 33390 32970
rect 33480 32910 33630 32970
rect 33480 32880 33540 32910
rect 34770 32880 34830 32970
rect 34920 32910 35070 32970
rect 34920 32880 34980 32910
rect 36210 32880 36270 32970
rect 36360 32910 36510 32970
rect 37650 32970 37710 33810
rect 37890 33090 37950 34320
rect 39090 33090 39150 34320
rect 37890 32970 37980 33090
rect 39060 32970 39150 33090
rect 39330 33930 39390 34320
rect 39330 33810 39420 33930
rect 39330 32970 39390 33810
rect 40680 34050 40740 34320
rect 40290 33570 40350 33720
rect 40440 33690 40500 33720
rect 40440 33630 40590 33690
rect 40200 33510 40350 33570
rect 40200 33090 40260 33510
rect 40530 33390 40590 33630
rect 40500 33270 40590 33390
rect 37650 32910 37800 32970
rect 36360 32880 36420 32910
rect 37740 32880 37800 32910
rect 37890 32880 37950 32970
rect 39090 32880 39150 32970
rect 39240 32910 39390 32970
rect 39240 32880 39300 32910
rect 40290 32880 40350 33030
rect 40530 32880 40590 33270
rect 40770 32880 40830 33990
rect 41730 33090 41790 34320
rect 41700 32970 41790 33090
rect 41970 33930 42030 34320
rect 41970 33810 42060 33930
rect 41970 32970 42030 33810
rect 43560 34050 43620 34320
rect 43170 33570 43230 33720
rect 43320 33690 43380 33720
rect 43320 33630 43470 33690
rect 43080 33510 43230 33570
rect 43080 33090 43140 33510
rect 43410 33390 43470 33630
rect 43380 33270 43470 33390
rect 41730 32880 41790 32970
rect 41880 32910 42030 32970
rect 41880 32880 41940 32910
rect 43170 32880 43230 33030
rect 43410 32880 43470 33270
rect 43650 32880 43710 33990
rect 46680 34050 46740 34320
rect 44370 33210 44430 33720
rect 44640 33690 44700 33720
rect 44610 33630 44700 33690
rect 44610 33510 44670 33630
rect 44370 32880 44430 33090
rect 44580 32970 44640 33390
rect 44790 33270 44850 33720
rect 45150 33540 45210 33720
rect 45300 33690 45360 33720
rect 45570 33690 45630 33720
rect 45300 33630 45630 33690
rect 45150 33480 45360 33540
rect 45300 33210 45360 33480
rect 45570 33210 45630 33630
rect 46290 33570 46350 33720
rect 46440 33690 46500 33720
rect 46440 33630 46590 33690
rect 46200 33510 46350 33570
rect 44880 33150 45120 33210
rect 44580 32910 44700 32970
rect 44640 32880 44700 32910
rect 44790 32910 44820 33030
rect 45060 32970 45120 33150
rect 46200 33090 46260 33510
rect 46530 33390 46590 33630
rect 46500 33270 46590 33390
rect 45570 32970 45630 33090
rect 45060 32910 45210 32970
rect 44790 32880 44850 32910
rect 45150 32880 45210 32910
rect 45300 32910 45630 32970
rect 45300 32880 45360 32910
rect 45570 32880 45630 32910
rect 46290 32880 46350 33030
rect 46530 32880 46590 33270
rect 46770 32880 46830 33990
rect 47730 33930 47790 34320
rect 47700 33810 47790 33930
rect 47730 32970 47790 33810
rect 47970 33090 48030 34320
rect 49170 33930 49230 34320
rect 49140 33810 49230 33930
rect 47970 32970 48060 33090
rect 49170 32970 49230 33810
rect 49410 33090 49470 34320
rect 49410 32970 49500 33090
rect 47730 32910 47880 32970
rect 47820 32880 47880 32910
rect 47970 32880 48030 32970
rect 49170 32910 49320 32970
rect 49260 32880 49320 32910
rect 49410 32880 49470 32970
rect 30450 32670 30540 32790
rect 30450 32580 30510 32670
rect 6690 32220 6750 32280
rect 6930 32220 6990 32280
rect 7170 32220 7230 32280
rect 7890 32220 7950 32280
rect 8130 32220 8190 32280
rect 8370 32220 8430 32280
rect 9090 32220 9150 32280
rect 9360 32220 9420 32280
rect 9510 32220 9570 32280
rect 9870 32220 9930 32280
rect 10020 32220 10080 32280
rect 10290 32220 10350 32280
rect 11250 32220 11310 32280
rect 11520 32220 11580 32280
rect 11670 32220 11730 32280
rect 12030 32220 12090 32280
rect 12180 32220 12240 32280
rect 12450 32220 12510 32280
rect 13890 32220 13950 32280
rect 15330 32220 15390 32280
rect 15480 32220 15540 32280
rect 16770 32220 16830 32280
rect 17010 32220 17070 32280
rect 17250 32220 17310 32280
rect 19500 32220 19560 32280
rect 19650 32220 19710 32280
rect 20940 32220 21000 32280
rect 21180 32220 21240 32280
rect 21330 32220 21390 32280
rect 23490 32220 23550 32280
rect 23730 32220 23790 32280
rect 23970 32220 24030 32280
rect 24930 32220 24990 32280
rect 25170 32220 25230 32280
rect 25410 32220 25470 32280
rect 26130 32220 26190 32280
rect 26400 32220 26460 32280
rect 26550 32220 26610 32280
rect 26910 32220 26970 32280
rect 27060 32220 27120 32280
rect 27330 32220 27390 32280
rect 30450 32220 30510 32280
rect 31260 32220 31320 32280
rect 31410 32220 31470 32280
rect 32130 32220 32190 32280
rect 32370 32220 32430 32280
rect 32610 32220 32670 32280
rect 33330 32220 33390 32280
rect 33480 32220 33540 32280
rect 34770 32220 34830 32280
rect 34920 32220 34980 32280
rect 36210 32220 36270 32280
rect 36360 32220 36420 32280
rect 37740 32220 37800 32280
rect 37890 32220 37950 32280
rect 39090 32220 39150 32280
rect 39240 32220 39300 32280
rect 40290 32220 40350 32280
rect 40530 32220 40590 32280
rect 40770 32220 40830 32280
rect 41730 32220 41790 32280
rect 41880 32220 41940 32280
rect 43170 32220 43230 32280
rect 43410 32220 43470 32280
rect 43650 32220 43710 32280
rect 44370 32220 44430 32280
rect 44640 32220 44700 32280
rect 44790 32220 44850 32280
rect 45150 32220 45210 32280
rect 45300 32220 45360 32280
rect 45570 32220 45630 32280
rect 46290 32220 46350 32280
rect 46530 32220 46590 32280
rect 46770 32220 46830 32280
rect 47820 32220 47880 32280
rect 47970 32220 48030 32280
rect 49260 32220 49320 32280
rect 49410 32220 49470 32280
rect 5490 31920 5550 31980
rect 5760 31920 5820 31980
rect 5910 31920 5970 31980
rect 6270 31920 6330 31980
rect 6420 31920 6480 31980
rect 6690 31920 6750 31980
rect 8130 31920 8190 31980
rect 8370 31920 8430 31980
rect 8610 31920 8670 31980
rect 9900 31920 9960 31980
rect 10050 31920 10110 31980
rect 11250 31920 11310 31980
rect 11520 31920 11580 31980
rect 11670 31920 11730 31980
rect 12030 31920 12090 31980
rect 12180 31920 12240 31980
rect 12450 31920 12510 31980
rect 14850 31920 14910 31980
rect 15120 31920 15180 31980
rect 15270 31920 15330 31980
rect 15630 31920 15690 31980
rect 15780 31920 15840 31980
rect 16050 31920 16110 31980
rect 17250 31920 17310 31980
rect 17520 31920 17580 31980
rect 17670 31920 17730 31980
rect 18030 31920 18090 31980
rect 18180 31920 18240 31980
rect 18450 31920 18510 31980
rect 19410 31920 19470 31980
rect 19680 31920 19740 31980
rect 19830 31920 19890 31980
rect 20190 31920 20250 31980
rect 20340 31920 20400 31980
rect 20610 31920 20670 31980
rect 21330 31920 21390 31980
rect 21480 31920 21540 31980
rect 22290 31920 22350 31980
rect 22530 31920 22590 31980
rect 22770 31920 22830 31980
rect 23970 31920 24030 31980
rect 25020 31920 25080 31980
rect 25260 31920 25320 31980
rect 25410 31920 25470 31980
rect 26130 31920 26190 31980
rect 26370 31920 26430 31980
rect 26610 31920 26670 31980
rect 27330 31920 27390 31980
rect 27900 31920 27960 31980
rect 28050 31920 28110 31980
rect 28770 31920 28830 31980
rect 29250 31920 29310 31980
rect 29490 31920 29550 31980
rect 29730 31920 29790 31980
rect 30930 31920 30990 31980
rect 31200 31920 31260 31980
rect 31350 31920 31410 31980
rect 31710 31920 31770 31980
rect 31860 31920 31920 31980
rect 32130 31920 32190 31980
rect 33330 31920 33390 31980
rect 33480 31920 33540 31980
rect 34770 31920 34830 31980
rect 34920 31920 34980 31980
rect 36210 31920 36270 31980
rect 36450 31920 36510 31980
rect 36690 31920 36750 31980
rect 37890 31920 37950 31980
rect 38040 31920 38100 31980
rect 39090 31920 39150 31980
rect 39330 31920 39390 31980
rect 39570 31920 39630 31980
rect 40770 31920 40830 31980
rect 41820 31920 41880 31980
rect 41970 31920 42030 31980
rect 43170 31920 43230 31980
rect 43410 31920 43470 31980
rect 43650 31920 43710 31980
rect 44610 31920 44670 31980
rect 44850 31920 44910 31980
rect 45090 31920 45150 31980
rect 46380 31920 46440 31980
rect 46530 31920 46590 31980
rect 48210 31920 48270 31980
rect 48480 31920 48540 31980
rect 48630 31920 48690 31980
rect 48990 31920 49050 31980
rect 49140 31920 49200 31980
rect 49410 31920 49470 31980
rect 23970 31530 24030 31620
rect 23970 31410 24060 31530
rect 5490 31290 5550 31320
rect 5760 31290 5820 31320
rect 5490 31230 5820 31290
rect 5910 31290 5970 31320
rect 6270 31290 6330 31320
rect 5910 31230 6060 31290
rect 5490 31110 5550 31230
rect 6000 31050 6060 31230
rect 6300 31230 6330 31290
rect 6420 31290 6480 31320
rect 6420 31230 6540 31290
rect 6000 30990 6210 31050
rect 5490 30570 5550 30990
rect 5820 30900 5880 30990
rect 5820 30840 5970 30900
rect 5490 30510 5820 30570
rect 5490 30480 5550 30510
rect 5760 30480 5820 30510
rect 5910 30480 5970 30840
rect 6150 30690 6210 30990
rect 6480 30870 6540 31230
rect 6690 31110 6750 31320
rect 8130 31170 8190 31320
rect 6270 30480 6330 30690
rect 6480 30570 6540 30750
rect 6720 30600 6780 30990
rect 8040 30690 8100 31110
rect 8370 30930 8430 31320
rect 8340 30810 8430 30930
rect 8040 30630 8190 30690
rect 6420 30510 6540 30570
rect 6690 30540 6780 30600
rect 6420 30480 6480 30510
rect 6690 30480 6750 30540
rect 8130 30480 8190 30630
rect 8370 30570 8430 30810
rect 8280 30510 8430 30570
rect 8280 30480 8340 30510
rect 8610 30210 8670 31320
rect 9900 31290 9960 31320
rect 9810 31230 9960 31290
rect 10050 31230 10110 31320
rect 9810 30390 9870 31230
rect 9780 30270 9870 30390
rect 8520 29880 8580 30150
rect 9810 29880 9870 30270
rect 10050 31110 10140 31230
rect 11250 31110 11310 31320
rect 11520 31290 11580 31320
rect 11460 31230 11580 31290
rect 11670 31290 11730 31320
rect 12030 31290 12090 31320
rect 10050 29880 10110 31110
rect 11250 30480 11310 30990
rect 11460 30810 11520 31230
rect 11670 31170 11700 31290
rect 11940 31230 12090 31290
rect 12180 31290 12240 31320
rect 12450 31290 12510 31320
rect 12180 31230 12510 31290
rect 11940 31050 12000 31230
rect 12450 31110 12510 31230
rect 14850 31110 14910 31320
rect 15120 31290 15180 31320
rect 15060 31230 15180 31290
rect 15270 31290 15330 31320
rect 15630 31290 15690 31320
rect 15270 31230 15300 31290
rect 11760 30990 12000 31050
rect 11490 30570 11550 30690
rect 11490 30510 11580 30570
rect 11520 30480 11580 30510
rect 11670 30480 11730 30930
rect 12180 30720 12240 30990
rect 12030 30660 12240 30720
rect 12030 30480 12090 30660
rect 12450 30570 12510 30990
rect 12180 30510 12510 30570
rect 14820 30600 14880 30990
rect 15060 30870 15120 31230
rect 15540 31230 15690 31290
rect 15780 31290 15840 31320
rect 16050 31290 16110 31320
rect 15780 31230 16110 31290
rect 15540 31050 15600 31230
rect 16050 31110 16110 31230
rect 17250 31110 17310 31320
rect 17520 31290 17580 31320
rect 17460 31230 17580 31290
rect 17670 31290 17730 31320
rect 18030 31290 18090 31320
rect 17670 31230 17700 31290
rect 14820 30540 14910 30600
rect 12180 30480 12240 30510
rect 12450 30480 12510 30510
rect 14850 30480 14910 30540
rect 15060 30570 15120 30750
rect 15390 30990 15600 31050
rect 15390 30690 15450 30990
rect 15720 30900 15780 30990
rect 15060 30510 15180 30570
rect 15120 30480 15180 30510
rect 15270 30480 15330 30690
rect 15630 30840 15780 30900
rect 15630 30480 15690 30840
rect 16050 30570 16110 30990
rect 15780 30510 16110 30570
rect 17220 30600 17280 30990
rect 17460 30870 17520 31230
rect 17940 31230 18090 31290
rect 18180 31290 18240 31320
rect 18450 31290 18510 31320
rect 18180 31230 18510 31290
rect 17940 31050 18000 31230
rect 18450 31110 18510 31230
rect 19410 31110 19470 31320
rect 19680 31290 19740 31320
rect 19620 31230 19740 31290
rect 19830 31290 19890 31320
rect 20190 31290 20250 31320
rect 17220 30540 17310 30600
rect 15780 30480 15840 30510
rect 16050 30480 16110 30510
rect 17250 30480 17310 30540
rect 17460 30570 17520 30750
rect 17790 30990 18000 31050
rect 17790 30690 17850 30990
rect 18120 30900 18180 30990
rect 17460 30510 17580 30570
rect 17520 30480 17580 30510
rect 17670 30480 17730 30690
rect 18030 30840 18180 30900
rect 18030 30480 18090 30840
rect 18450 30570 18510 30990
rect 18180 30510 18510 30570
rect 18180 30480 18240 30510
rect 18450 30480 18510 30510
rect 19410 30480 19470 30990
rect 19620 30810 19680 31230
rect 19830 31170 19860 31290
rect 20100 31230 20250 31290
rect 20340 31290 20400 31320
rect 20610 31290 20670 31320
rect 20340 31230 20670 31290
rect 21330 31230 21390 31320
rect 21480 31290 21540 31320
rect 21480 31230 21630 31290
rect 20100 31050 20160 31230
rect 20610 31110 20670 31230
rect 21300 31110 21390 31230
rect 19920 30990 20160 31050
rect 19650 30570 19710 30690
rect 19650 30510 19740 30570
rect 19680 30480 19740 30510
rect 19830 30480 19890 30930
rect 20340 30720 20400 30990
rect 20190 30660 20400 30720
rect 20190 30480 20250 30660
rect 20610 30570 20670 30990
rect 20340 30510 20670 30570
rect 20340 30480 20400 30510
rect 20610 30480 20670 30510
rect 21330 29880 21390 31110
rect 21570 30390 21630 31230
rect 21570 30270 21660 30390
rect 21570 29880 21630 30270
rect 22290 30210 22350 31320
rect 22530 30930 22590 31320
rect 22770 31170 22830 31320
rect 22530 30810 22620 30930
rect 22530 30570 22590 30810
rect 22860 30690 22920 31110
rect 22770 30630 22920 30690
rect 22530 30510 22680 30570
rect 22620 30480 22680 30510
rect 22770 30480 22830 30630
rect 22380 29880 22440 30150
rect 23970 29880 24030 31410
rect 25020 31230 25080 31620
rect 27330 31530 27390 31620
rect 27330 31410 27420 31530
rect 24930 31110 24960 31200
rect 24930 29880 24990 31110
rect 25260 30990 25320 31320
rect 25170 30930 25320 30990
rect 25410 30990 25470 31320
rect 25170 30630 25230 30930
rect 25410 30870 25500 30990
rect 25170 29880 25230 30510
rect 25410 29880 25470 30870
rect 26130 30210 26190 31320
rect 26370 30930 26430 31320
rect 26610 31170 26670 31320
rect 26370 30810 26460 30930
rect 26370 30570 26430 30810
rect 26700 30690 26760 31110
rect 26610 30630 26760 30690
rect 26370 30510 26520 30570
rect 26460 30480 26520 30510
rect 26610 30480 26670 30630
rect 26220 29880 26280 30150
rect 27330 29880 27390 31410
rect 28770 31530 28830 31620
rect 28740 31410 28830 31530
rect 27900 31290 27960 31320
rect 27810 31230 27960 31290
rect 28050 31230 28110 31320
rect 27810 30390 27870 31230
rect 27780 30270 27870 30390
rect 27810 29880 27870 30270
rect 28050 31110 28140 31230
rect 28050 29880 28110 31110
rect 28770 29880 28830 31410
rect 40770 31530 40830 31620
rect 40770 31410 40860 31530
rect 29250 30210 29310 31320
rect 29490 30930 29550 31320
rect 29730 31170 29790 31320
rect 30930 31290 30990 31320
rect 31200 31290 31260 31320
rect 30930 31230 31260 31290
rect 31350 31290 31410 31320
rect 31710 31290 31770 31320
rect 31350 31230 31500 31290
rect 30930 31110 30990 31230
rect 29490 30810 29580 30930
rect 29490 30570 29550 30810
rect 29820 30690 29880 31110
rect 31440 31050 31500 31230
rect 31740 31170 31770 31290
rect 31860 31290 31920 31320
rect 31860 31230 31980 31290
rect 31440 30990 31680 31050
rect 29730 30630 29880 30690
rect 29490 30510 29640 30570
rect 29580 30480 29640 30510
rect 29730 30480 29790 30630
rect 30930 30570 30990 30990
rect 31200 30720 31260 30990
rect 31200 30660 31410 30720
rect 30930 30510 31260 30570
rect 30930 30480 30990 30510
rect 31200 30480 31260 30510
rect 31350 30480 31410 30660
rect 31710 30480 31770 30930
rect 31920 30810 31980 31230
rect 32130 31110 32190 31320
rect 33330 31230 33390 31320
rect 33480 31290 33540 31320
rect 33480 31230 33630 31290
rect 34770 31230 34830 31320
rect 34920 31290 34980 31320
rect 34920 31230 35070 31290
rect 33300 31110 33390 31230
rect 31890 30570 31950 30690
rect 31860 30510 31950 30570
rect 31860 30480 31920 30510
rect 32130 30480 32190 30990
rect 29340 29880 29400 30150
rect 33330 29880 33390 31110
rect 33570 30390 33630 31230
rect 34740 31110 34830 31230
rect 33570 30270 33660 30390
rect 33570 29880 33630 30270
rect 34770 29880 34830 31110
rect 35010 30390 35070 31230
rect 35010 30270 35100 30390
rect 35010 29880 35070 30270
rect 36210 30210 36270 31320
rect 36450 30930 36510 31320
rect 36690 31170 36750 31320
rect 37890 31230 37950 31320
rect 38040 31290 38100 31320
rect 38040 31230 38190 31290
rect 37860 31110 37950 31230
rect 36450 30810 36540 30930
rect 36450 30570 36510 30810
rect 36780 30690 36840 31110
rect 36690 30630 36840 30690
rect 36450 30510 36600 30570
rect 36540 30480 36600 30510
rect 36690 30480 36750 30630
rect 36300 29880 36360 30150
rect 37890 29880 37950 31110
rect 38130 30390 38190 31230
rect 39090 31170 39150 31320
rect 39000 30690 39060 31110
rect 39330 30930 39390 31320
rect 39300 30810 39390 30930
rect 39000 30630 39150 30690
rect 39090 30480 39150 30630
rect 39330 30570 39390 30810
rect 39240 30510 39390 30570
rect 39240 30480 39300 30510
rect 38130 30270 38220 30390
rect 38130 29880 38190 30270
rect 39570 30210 39630 31320
rect 39480 29880 39540 30150
rect 40770 29880 40830 31410
rect 41820 31290 41880 31320
rect 41730 31230 41880 31290
rect 41970 31230 42030 31320
rect 41730 30390 41790 31230
rect 41700 30270 41790 30390
rect 41730 29880 41790 30270
rect 41970 31110 42060 31230
rect 41970 29880 42030 31110
rect 43170 30210 43230 31320
rect 43410 30930 43470 31320
rect 43650 31170 43710 31320
rect 44610 31170 44670 31320
rect 43410 30810 43500 30930
rect 43410 30570 43470 30810
rect 43740 30690 43800 31110
rect 43650 30630 43800 30690
rect 44520 30690 44580 31110
rect 44850 30930 44910 31320
rect 44820 30810 44910 30930
rect 44520 30630 44670 30690
rect 43410 30510 43560 30570
rect 43500 30480 43560 30510
rect 43650 30480 43710 30630
rect 44610 30480 44670 30630
rect 44850 30570 44910 30810
rect 44760 30510 44910 30570
rect 44760 30480 44820 30510
rect 43260 29880 43320 30150
rect 45090 30210 45150 31320
rect 46380 31290 46440 31320
rect 46290 31230 46440 31290
rect 46530 31230 46590 31320
rect 46290 30390 46350 31230
rect 46260 30270 46350 30390
rect 45000 29880 45060 30150
rect 46290 29880 46350 30270
rect 46530 31110 46620 31230
rect 48210 31110 48270 31320
rect 48480 31290 48540 31320
rect 48420 31230 48540 31290
rect 48630 31290 48690 31320
rect 48990 31290 49050 31320
rect 46530 29880 46590 31110
rect 48210 30480 48270 30990
rect 48420 30810 48480 31230
rect 48630 31170 48660 31290
rect 48900 31230 49050 31290
rect 49140 31290 49200 31320
rect 49410 31290 49470 31320
rect 49140 31230 49470 31290
rect 48900 31050 48960 31230
rect 49410 31110 49470 31230
rect 48720 30990 48960 31050
rect 48450 30570 48510 30690
rect 48450 30510 48540 30570
rect 48480 30480 48540 30510
rect 48630 30480 48690 30930
rect 49140 30720 49200 30990
rect 48990 30660 49200 30720
rect 48990 30480 49050 30660
rect 49410 30570 49470 30990
rect 49140 30510 49470 30570
rect 49140 30480 49200 30510
rect 49410 30480 49470 30510
rect 5490 29220 5550 29280
rect 5760 29220 5820 29280
rect 5910 29220 5970 29280
rect 6270 29220 6330 29280
rect 6420 29220 6480 29280
rect 6690 29220 6750 29280
rect 8130 29220 8190 29280
rect 8280 29220 8340 29280
rect 8520 29220 8580 29280
rect 9810 29220 9870 29280
rect 10050 29220 10110 29280
rect 11250 29220 11310 29280
rect 11520 29220 11580 29280
rect 11670 29220 11730 29280
rect 12030 29220 12090 29280
rect 12180 29220 12240 29280
rect 12450 29220 12510 29280
rect 14850 29220 14910 29280
rect 15120 29220 15180 29280
rect 15270 29220 15330 29280
rect 15630 29220 15690 29280
rect 15780 29220 15840 29280
rect 16050 29220 16110 29280
rect 17250 29220 17310 29280
rect 17520 29220 17580 29280
rect 17670 29220 17730 29280
rect 18030 29220 18090 29280
rect 18180 29220 18240 29280
rect 18450 29220 18510 29280
rect 19410 29220 19470 29280
rect 19680 29220 19740 29280
rect 19830 29220 19890 29280
rect 20190 29220 20250 29280
rect 20340 29220 20400 29280
rect 20610 29220 20670 29280
rect 21330 29220 21390 29280
rect 21570 29220 21630 29280
rect 22380 29220 22440 29280
rect 22620 29220 22680 29280
rect 22770 29220 22830 29280
rect 23970 29220 24030 29280
rect 24930 29220 24990 29280
rect 25170 29220 25230 29280
rect 25410 29220 25470 29280
rect 26220 29220 26280 29280
rect 26460 29220 26520 29280
rect 26610 29220 26670 29280
rect 27330 29220 27390 29280
rect 27810 29220 27870 29280
rect 28050 29220 28110 29280
rect 28770 29220 28830 29280
rect 29340 29220 29400 29280
rect 29580 29220 29640 29280
rect 29730 29220 29790 29280
rect 30930 29220 30990 29280
rect 31200 29220 31260 29280
rect 31350 29220 31410 29280
rect 31710 29220 31770 29280
rect 31860 29220 31920 29280
rect 32130 29220 32190 29280
rect 33330 29220 33390 29280
rect 33570 29220 33630 29280
rect 34770 29220 34830 29280
rect 35010 29220 35070 29280
rect 36300 29220 36360 29280
rect 36540 29220 36600 29280
rect 36690 29220 36750 29280
rect 37890 29220 37950 29280
rect 38130 29220 38190 29280
rect 39090 29220 39150 29280
rect 39240 29220 39300 29280
rect 39480 29220 39540 29280
rect 40770 29220 40830 29280
rect 41730 29220 41790 29280
rect 41970 29220 42030 29280
rect 43260 29220 43320 29280
rect 43500 29220 43560 29280
rect 43650 29220 43710 29280
rect 44610 29220 44670 29280
rect 44760 29220 44820 29280
rect 45000 29220 45060 29280
rect 46290 29220 46350 29280
rect 46530 29220 46590 29280
rect 48210 29220 48270 29280
rect 48480 29220 48540 29280
rect 48630 29220 48690 29280
rect 48990 29220 49050 29280
rect 49140 29220 49200 29280
rect 49410 29220 49470 29280
rect 7170 28920 7230 28980
rect 7440 28920 7500 28980
rect 7590 28920 7650 28980
rect 7950 28920 8010 28980
rect 8100 28920 8160 28980
rect 8370 28920 8430 28980
rect 8850 28920 8910 28980
rect 9090 28920 9150 28980
rect 9570 28920 9630 28980
rect 9840 28920 9900 28980
rect 9990 28920 10050 28980
rect 10350 28920 10410 28980
rect 10500 28920 10560 28980
rect 10770 28920 10830 28980
rect 11250 28920 11310 28980
rect 11400 28920 11460 28980
rect 11640 28920 11700 28980
rect 12210 28920 12270 28980
rect 12450 28920 12510 28980
rect 12930 28920 12990 28980
rect 13170 28920 13230 28980
rect 13890 28920 13950 28980
rect 14130 28920 14190 28980
rect 14370 28920 14430 28980
rect 15570 28920 15630 28980
rect 15810 28920 15870 28980
rect 16770 28920 16830 28980
rect 17010 28920 17070 28980
rect 18210 28920 18270 28980
rect 18450 28920 18510 28980
rect 19500 28920 19560 28980
rect 19740 28920 19800 28980
rect 19890 28920 19950 28980
rect 21090 28920 21150 28980
rect 21330 28920 21390 28980
rect 22290 28920 22350 28980
rect 22530 28920 22590 28980
rect 23730 28920 23790 28980
rect 23970 28920 24030 28980
rect 25170 28920 25230 28980
rect 25410 28920 25470 28980
rect 26610 28920 26670 28980
rect 26850 28920 26910 28980
rect 28620 28920 28680 28980
rect 28860 28920 28920 28980
rect 29010 28920 29070 28980
rect 30450 28920 30510 28980
rect 30690 28920 30750 28980
rect 31980 28920 32040 28980
rect 32220 28920 32280 28980
rect 32370 28920 32430 28980
rect 33090 28920 33150 28980
rect 33360 28920 33420 28980
rect 33510 28920 33570 28980
rect 33870 28920 33930 28980
rect 34020 28920 34080 28980
rect 34290 28920 34350 28980
rect 35010 28920 35070 28980
rect 35250 28920 35310 28980
rect 36210 28920 36270 28980
rect 36450 28920 36510 28980
rect 37650 28920 37710 28980
rect 37890 28920 37950 28980
rect 38850 28920 38910 28980
rect 39090 28920 39150 28980
rect 39810 28920 39870 28980
rect 40080 28920 40140 28980
rect 40230 28920 40290 28980
rect 40590 28920 40650 28980
rect 40740 28920 40800 28980
rect 41010 28920 41070 28980
rect 41730 28920 41790 28980
rect 41970 28920 42030 28980
rect 43260 28920 43320 28980
rect 43500 28920 43560 28980
rect 43650 28920 43710 28980
rect 44610 28920 44670 28980
rect 44760 28920 44820 28980
rect 45000 28920 45060 28980
rect 46050 28920 46110 28980
rect 46200 28920 46260 28980
rect 46440 28920 46500 28980
rect 47010 28920 47070 28980
rect 47490 28920 47550 28980
rect 47730 28920 47790 28980
rect 47970 28920 48030 28980
rect 48210 28920 48270 28980
rect 48690 28920 48750 28980
rect 48930 28920 48990 28980
rect 49410 28920 49470 28980
rect 49560 28920 49620 28980
rect 49800 28920 49860 28980
rect 7170 27210 7230 27720
rect 7440 27690 7500 27720
rect 7410 27630 7500 27690
rect 7410 27510 7470 27630
rect 7170 26880 7230 27090
rect 7380 26970 7440 27390
rect 7590 27270 7650 27720
rect 7950 27540 8010 27720
rect 8100 27690 8160 27720
rect 8370 27690 8430 27720
rect 8100 27630 8430 27690
rect 7950 27480 8160 27540
rect 8100 27210 8160 27480
rect 8370 27210 8430 27630
rect 7680 27150 7920 27210
rect 7380 26910 7500 26970
rect 7440 26880 7500 26910
rect 7590 26910 7620 27030
rect 7860 26970 7920 27150
rect 8850 27090 8910 28320
rect 8370 26970 8430 27090
rect 8820 26970 8910 27090
rect 9090 27930 9150 28320
rect 9090 27810 9180 27930
rect 9090 26970 9150 27810
rect 11640 28050 11700 28320
rect 9570 27690 9630 27720
rect 9840 27690 9900 27720
rect 9570 27630 9900 27690
rect 9570 27210 9630 27630
rect 9990 27360 10050 27720
rect 9900 27300 10050 27360
rect 10350 27510 10410 27720
rect 10500 27690 10560 27720
rect 10500 27630 10620 27690
rect 9900 27210 9960 27300
rect 10230 27210 10290 27510
rect 10080 27150 10290 27210
rect 10560 27450 10620 27630
rect 10770 27660 10830 27720
rect 10770 27600 10860 27660
rect 7860 26910 8010 26970
rect 7590 26880 7650 26910
rect 7950 26880 8010 26910
rect 8100 26910 8430 26970
rect 8100 26880 8160 26910
rect 8370 26880 8430 26910
rect 8850 26880 8910 26970
rect 9000 26910 9150 26970
rect 9570 26970 9630 27090
rect 10080 26970 10140 27150
rect 9570 26910 9900 26970
rect 9000 26880 9060 26910
rect 9570 26880 9630 26910
rect 9840 26880 9900 26910
rect 9990 26910 10140 26970
rect 10560 26970 10620 27330
rect 10800 27210 10860 27600
rect 11250 27570 11310 27720
rect 11400 27690 11460 27720
rect 11400 27630 11550 27690
rect 11160 27510 11310 27570
rect 11160 27090 11220 27510
rect 11490 27390 11550 27630
rect 11460 27270 11550 27390
rect 10380 26910 10410 26970
rect 9990 26880 10050 26910
rect 10350 26880 10410 26910
rect 10500 26910 10620 26970
rect 10500 26880 10560 26910
rect 10770 26880 10830 27090
rect 11250 26880 11310 27030
rect 11490 26880 11550 27270
rect 11730 26880 11790 27990
rect 12210 27090 12270 28320
rect 12180 26970 12270 27090
rect 12450 27930 12510 28320
rect 12450 27810 12540 27930
rect 12450 26970 12510 27810
rect 12930 27090 12990 28320
rect 12900 26970 12990 27090
rect 13170 27930 13230 28320
rect 13170 27810 13260 27930
rect 13170 26970 13230 27810
rect 13890 27090 13950 28320
rect 14130 27690 14190 28320
rect 14130 27270 14190 27570
rect 14370 27330 14430 28320
rect 14130 27210 14280 27270
rect 13890 27000 13920 27090
rect 12210 26880 12270 26970
rect 12360 26910 12510 26970
rect 12360 26880 12420 26910
rect 12930 26880 12990 26970
rect 13080 26910 13230 26970
rect 13080 26880 13140 26910
rect 13980 26580 14040 26970
rect 14220 26880 14280 27210
rect 14370 27210 14460 27330
rect 14370 26880 14430 27210
rect 15570 27090 15630 28320
rect 15540 26970 15630 27090
rect 15810 27930 15870 28320
rect 16770 27930 16830 28320
rect 15810 27810 15900 27930
rect 16740 27810 16830 27930
rect 15810 26970 15870 27810
rect 15570 26880 15630 26970
rect 15720 26910 15870 26970
rect 16770 26970 16830 27810
rect 17010 27090 17070 28320
rect 18210 27090 18270 28320
rect 17010 26970 17100 27090
rect 18180 26970 18270 27090
rect 18450 27930 18510 28320
rect 19500 28050 19560 28320
rect 18450 27810 18540 27930
rect 18450 26970 18510 27810
rect 16770 26910 16920 26970
rect 15720 26880 15780 26910
rect 16860 26880 16920 26910
rect 17010 26880 17070 26970
rect 18210 26880 18270 26970
rect 18360 26910 18510 26970
rect 18360 26880 18420 26910
rect 19410 26880 19470 27990
rect 19740 27690 19800 27720
rect 19650 27630 19800 27690
rect 19650 27390 19710 27630
rect 19890 27570 19950 27720
rect 19890 27510 20040 27570
rect 19650 27270 19740 27390
rect 19650 26880 19710 27270
rect 19980 27090 20040 27510
rect 21090 27090 21150 28320
rect 19890 26880 19950 27030
rect 21060 26970 21150 27090
rect 21330 27930 21390 28320
rect 21330 27810 21420 27930
rect 21330 26970 21390 27810
rect 22290 27090 22350 28320
rect 22260 26970 22350 27090
rect 22530 27930 22590 28320
rect 22530 27810 22620 27930
rect 22530 26970 22590 27810
rect 23730 27090 23790 28320
rect 23700 26970 23790 27090
rect 23970 27930 24030 28320
rect 23970 27810 24060 27930
rect 23970 26970 24030 27810
rect 25170 27090 25230 28320
rect 25140 26970 25230 27090
rect 25410 27930 25470 28320
rect 25410 27810 25500 27930
rect 25410 26970 25470 27810
rect 26610 27090 26670 28320
rect 26580 26970 26670 27090
rect 26850 27930 26910 28320
rect 28620 28050 28680 28320
rect 26850 27810 26940 27930
rect 26850 26970 26910 27810
rect 21090 26880 21150 26970
rect 21240 26910 21390 26970
rect 21240 26880 21300 26910
rect 22290 26880 22350 26970
rect 22440 26910 22590 26970
rect 22440 26880 22500 26910
rect 23730 26880 23790 26970
rect 23880 26910 24030 26970
rect 23880 26880 23940 26910
rect 25170 26880 25230 26970
rect 25320 26910 25470 26970
rect 25320 26880 25380 26910
rect 26610 26880 26670 26970
rect 26760 26910 26910 26970
rect 26760 26880 26820 26910
rect 28530 26880 28590 27990
rect 30450 27930 30510 28320
rect 30420 27810 30510 27930
rect 28860 27690 28920 27720
rect 28770 27630 28920 27690
rect 28770 27390 28830 27630
rect 29010 27570 29070 27720
rect 29010 27510 29160 27570
rect 28770 27270 28860 27390
rect 28770 26880 28830 27270
rect 29100 27090 29160 27510
rect 29010 26880 29070 27030
rect 30450 26970 30510 27810
rect 30690 27090 30750 28320
rect 31980 28050 32040 28320
rect 30690 26970 30780 27090
rect 30450 26910 30600 26970
rect 30540 26880 30600 26910
rect 30690 26880 30750 26970
rect 31890 26880 31950 27990
rect 32220 27690 32280 27720
rect 32130 27630 32280 27690
rect 32130 27390 32190 27630
rect 32370 27570 32430 27720
rect 32370 27510 32520 27570
rect 32130 27270 32220 27390
rect 32130 26880 32190 27270
rect 32460 27090 32520 27510
rect 33090 27210 33150 27720
rect 33360 27690 33420 27720
rect 33330 27630 33420 27690
rect 33330 27510 33390 27630
rect 32370 26880 32430 27030
rect 33090 26880 33150 27090
rect 33300 26970 33360 27390
rect 33510 27270 33570 27720
rect 33870 27540 33930 27720
rect 34020 27690 34080 27720
rect 34290 27690 34350 27720
rect 34020 27630 34350 27690
rect 33870 27480 34080 27540
rect 34020 27210 34080 27480
rect 34290 27210 34350 27630
rect 33600 27150 33840 27210
rect 33300 26910 33420 26970
rect 33360 26880 33420 26910
rect 33510 26910 33540 27030
rect 33780 26970 33840 27150
rect 35010 27090 35070 28320
rect 34290 26970 34350 27090
rect 34980 26970 35070 27090
rect 35250 27930 35310 28320
rect 35250 27810 35340 27930
rect 35250 26970 35310 27810
rect 36210 27090 36270 28320
rect 36180 26970 36270 27090
rect 36450 27930 36510 28320
rect 37650 27930 37710 28320
rect 36450 27810 36540 27930
rect 37620 27810 37710 27930
rect 36450 26970 36510 27810
rect 33780 26910 33930 26970
rect 33510 26880 33570 26910
rect 33870 26880 33930 26910
rect 34020 26910 34350 26970
rect 34020 26880 34080 26910
rect 34290 26880 34350 26910
rect 35010 26880 35070 26970
rect 35160 26910 35310 26970
rect 35160 26880 35220 26910
rect 36210 26880 36270 26970
rect 36360 26910 36510 26970
rect 37650 26970 37710 27810
rect 37890 27090 37950 28320
rect 38850 27090 38910 28320
rect 37890 26970 37980 27090
rect 38820 26970 38910 27090
rect 39090 27930 39150 28320
rect 39090 27810 39180 27930
rect 39090 26970 39150 27810
rect 39810 27210 39870 27720
rect 40080 27690 40140 27720
rect 40050 27630 40140 27690
rect 40050 27510 40110 27630
rect 37650 26910 37800 26970
rect 36360 26880 36420 26910
rect 37740 26880 37800 26910
rect 37890 26880 37950 26970
rect 38850 26880 38910 26970
rect 39000 26910 39150 26970
rect 39000 26880 39060 26910
rect 39810 26880 39870 27090
rect 40020 26970 40080 27390
rect 40230 27270 40290 27720
rect 40590 27540 40650 27720
rect 40740 27690 40800 27720
rect 41010 27690 41070 27720
rect 40740 27630 41070 27690
rect 40590 27480 40800 27540
rect 40740 27210 40800 27480
rect 41010 27210 41070 27630
rect 40320 27150 40560 27210
rect 40020 26910 40140 26970
rect 40080 26880 40140 26910
rect 40230 26910 40260 27030
rect 40500 26970 40560 27150
rect 41730 27090 41790 28320
rect 41010 26970 41070 27090
rect 41700 26970 41790 27090
rect 41970 27930 42030 28320
rect 43260 28050 43320 28320
rect 41970 27810 42060 27930
rect 41970 26970 42030 27810
rect 40500 26910 40650 26970
rect 40230 26880 40290 26910
rect 40590 26880 40650 26910
rect 40740 26910 41070 26970
rect 40740 26880 40800 26910
rect 41010 26880 41070 26910
rect 41730 26880 41790 26970
rect 41880 26910 42030 26970
rect 41880 26880 41940 26910
rect 43170 26880 43230 27990
rect 45000 28050 45060 28320
rect 43500 27690 43560 27720
rect 43410 27630 43560 27690
rect 43410 27390 43470 27630
rect 43650 27570 43710 27720
rect 44610 27570 44670 27720
rect 44760 27690 44820 27720
rect 44760 27630 44910 27690
rect 43650 27510 43800 27570
rect 43410 27270 43500 27390
rect 43410 26880 43470 27270
rect 43740 27090 43800 27510
rect 44520 27510 44670 27570
rect 44520 27090 44580 27510
rect 44850 27390 44910 27630
rect 44820 27270 44910 27390
rect 43650 26880 43710 27030
rect 44610 26880 44670 27030
rect 44850 26880 44910 27270
rect 45090 26880 45150 27990
rect 46440 28050 46500 28320
rect 46050 27570 46110 27720
rect 46200 27690 46260 27720
rect 46200 27630 46350 27690
rect 45960 27510 46110 27570
rect 45960 27090 46020 27510
rect 46290 27390 46350 27630
rect 46260 27270 46350 27390
rect 46050 26880 46110 27030
rect 46290 26880 46350 27270
rect 46530 26880 46590 27990
rect 47010 26790 47070 28320
rect 47490 27690 47550 27720
rect 47430 27630 47550 27690
rect 47460 27510 47490 27630
rect 47430 27030 47490 27510
rect 47730 27300 47790 27720
rect 47970 27690 48030 27720
rect 47970 27630 48060 27690
rect 47730 27270 47760 27300
rect 47430 26970 47550 27030
rect 47700 26970 47760 27270
rect 47490 26880 47550 26970
rect 47640 26910 47760 26970
rect 47640 26880 47700 26910
rect 48000 26880 48060 27630
rect 48210 27570 48270 27720
rect 48300 26970 48360 27510
rect 48690 27090 48750 28320
rect 48660 26970 48750 27090
rect 48930 27930 48990 28320
rect 48930 27810 49020 27930
rect 48930 26970 48990 27810
rect 49800 28050 49860 28320
rect 49410 27570 49470 27720
rect 49560 27690 49620 27720
rect 49560 27630 49710 27690
rect 49320 27510 49470 27570
rect 49320 27090 49380 27510
rect 49650 27390 49710 27630
rect 49620 27270 49710 27390
rect 48150 26910 48360 26970
rect 48150 26880 48210 26910
rect 48690 26880 48750 26970
rect 48840 26910 48990 26970
rect 48840 26880 48900 26910
rect 49410 26880 49470 27030
rect 49650 26880 49710 27270
rect 49890 26880 49950 27990
rect 46980 26670 47070 26790
rect 47010 26580 47070 26670
rect 7170 26220 7230 26280
rect 7440 26220 7500 26280
rect 7590 26220 7650 26280
rect 7950 26220 8010 26280
rect 8100 26220 8160 26280
rect 8370 26220 8430 26280
rect 8850 26220 8910 26280
rect 9000 26220 9060 26280
rect 9570 26220 9630 26280
rect 9840 26220 9900 26280
rect 9990 26220 10050 26280
rect 10350 26220 10410 26280
rect 10500 26220 10560 26280
rect 10770 26220 10830 26280
rect 11250 26220 11310 26280
rect 11490 26220 11550 26280
rect 11730 26220 11790 26280
rect 12210 26220 12270 26280
rect 12360 26220 12420 26280
rect 12930 26220 12990 26280
rect 13080 26220 13140 26280
rect 13980 26220 14040 26280
rect 14220 26220 14280 26280
rect 14370 26220 14430 26280
rect 15570 26220 15630 26280
rect 15720 26220 15780 26280
rect 16860 26220 16920 26280
rect 17010 26220 17070 26280
rect 18210 26220 18270 26280
rect 18360 26220 18420 26280
rect 19410 26220 19470 26280
rect 19650 26220 19710 26280
rect 19890 26220 19950 26280
rect 21090 26220 21150 26280
rect 21240 26220 21300 26280
rect 22290 26220 22350 26280
rect 22440 26220 22500 26280
rect 23730 26220 23790 26280
rect 23880 26220 23940 26280
rect 25170 26220 25230 26280
rect 25320 26220 25380 26280
rect 26610 26220 26670 26280
rect 26760 26220 26820 26280
rect 28530 26220 28590 26280
rect 28770 26220 28830 26280
rect 29010 26220 29070 26280
rect 30540 26220 30600 26280
rect 30690 26220 30750 26280
rect 31890 26220 31950 26280
rect 32130 26220 32190 26280
rect 32370 26220 32430 26280
rect 33090 26220 33150 26280
rect 33360 26220 33420 26280
rect 33510 26220 33570 26280
rect 33870 26220 33930 26280
rect 34020 26220 34080 26280
rect 34290 26220 34350 26280
rect 35010 26220 35070 26280
rect 35160 26220 35220 26280
rect 36210 26220 36270 26280
rect 36360 26220 36420 26280
rect 37740 26220 37800 26280
rect 37890 26220 37950 26280
rect 38850 26220 38910 26280
rect 39000 26220 39060 26280
rect 39810 26220 39870 26280
rect 40080 26220 40140 26280
rect 40230 26220 40290 26280
rect 40590 26220 40650 26280
rect 40740 26220 40800 26280
rect 41010 26220 41070 26280
rect 41730 26220 41790 26280
rect 41880 26220 41940 26280
rect 43170 26220 43230 26280
rect 43410 26220 43470 26280
rect 43650 26220 43710 26280
rect 44610 26220 44670 26280
rect 44850 26220 44910 26280
rect 45090 26220 45150 26280
rect 46050 26220 46110 26280
rect 46290 26220 46350 26280
rect 46530 26220 46590 26280
rect 47010 26220 47070 26280
rect 47490 26220 47550 26280
rect 47640 26220 47700 26280
rect 48000 26220 48060 26280
rect 48150 26220 48210 26280
rect 48690 26220 48750 26280
rect 48840 26220 48900 26280
rect 49410 26220 49470 26280
rect 49650 26220 49710 26280
rect 49890 26220 49950 26280
rect 5490 25920 5550 25980
rect 5760 25920 5820 25980
rect 5910 25920 5970 25980
rect 6270 25920 6330 25980
rect 6420 25920 6480 25980
rect 6690 25920 6750 25980
rect 7170 25920 7230 25980
rect 7320 25920 7380 25980
rect 7890 25920 7950 25980
rect 8130 25920 8190 25980
rect 8370 25920 8430 25980
rect 8850 25920 8910 25980
rect 9000 25920 9060 25980
rect 9570 25920 9630 25980
rect 9840 25920 9900 25980
rect 9990 25920 10050 25980
rect 10350 25920 10410 25980
rect 10500 25920 10560 25980
rect 10770 25920 10830 25980
rect 12210 25920 12270 25980
rect 12450 25920 12510 25980
rect 12600 25920 12660 25980
rect 13890 25920 13950 25980
rect 15090 25920 15150 25980
rect 15330 25920 15390 25980
rect 15570 25920 15630 25980
rect 20940 25920 21000 25980
rect 21090 25920 21150 25980
rect 23250 25920 23310 25980
rect 23400 25920 23460 25980
rect 25650 25920 25710 25980
rect 25920 25920 25980 25980
rect 26070 25920 26130 25980
rect 26430 25920 26490 25980
rect 26580 25920 26640 25980
rect 26850 25920 26910 25980
rect 28050 25920 28110 25980
rect 28290 25920 28350 25980
rect 28530 25920 28590 25980
rect 30450 25920 30510 25980
rect 31170 25920 31230 25980
rect 31410 25920 31470 25980
rect 31650 25920 31710 25980
rect 32370 25920 32430 25980
rect 33330 25920 33390 25980
rect 33480 25920 33540 25980
rect 34770 25920 34830 25980
rect 34920 25920 34980 25980
rect 36210 25920 36270 25980
rect 36360 25920 36420 25980
rect 37650 25920 37710 25980
rect 37800 25920 37860 25980
rect 39090 25920 39150 25980
rect 39240 25920 39300 25980
rect 40530 25920 40590 25980
rect 40680 25920 40740 25980
rect 41970 25920 42030 25980
rect 42120 25920 42180 25980
rect 43410 25920 43470 25980
rect 43650 25920 43710 25980
rect 44610 25920 44670 25980
rect 47970 25920 48030 25980
rect 48240 25920 48300 25980
rect 48390 25920 48450 25980
rect 48750 25920 48810 25980
rect 48900 25920 48960 25980
rect 49170 25920 49230 25980
rect 5490 25110 5550 25320
rect 5760 25290 5820 25320
rect 5700 25230 5820 25290
rect 5910 25290 5970 25320
rect 6270 25290 6330 25320
rect 5490 24480 5550 24990
rect 5700 24810 5760 25230
rect 5910 25170 5940 25290
rect 6180 25230 6330 25290
rect 6420 25290 6480 25320
rect 6690 25290 6750 25320
rect 6420 25230 6750 25290
rect 7170 25230 7230 25320
rect 7320 25290 7380 25320
rect 7320 25230 7470 25290
rect 6180 25050 6240 25230
rect 6690 25110 6750 25230
rect 7140 25110 7230 25230
rect 6000 24990 6240 25050
rect 5730 24570 5790 24690
rect 5730 24510 5820 24570
rect 5760 24480 5820 24510
rect 5910 24480 5970 24930
rect 6420 24720 6480 24990
rect 6270 24660 6480 24720
rect 6270 24480 6330 24660
rect 6690 24570 6750 24990
rect 6420 24510 6750 24570
rect 6420 24480 6480 24510
rect 6690 24480 6750 24510
rect 7170 23880 7230 25110
rect 7410 24390 7470 25230
rect 7410 24270 7500 24390
rect 7410 23880 7470 24270
rect 7890 24210 7950 25320
rect 8130 24930 8190 25320
rect 8370 25170 8430 25320
rect 8850 25230 8910 25320
rect 9000 25290 9060 25320
rect 9000 25230 9150 25290
rect 8820 25110 8910 25230
rect 8130 24810 8220 24930
rect 8130 24570 8190 24810
rect 8460 24690 8520 25110
rect 8370 24630 8520 24690
rect 8130 24510 8280 24570
rect 8220 24480 8280 24510
rect 8370 24480 8430 24630
rect 7980 23880 8040 24150
rect 8850 23880 8910 25110
rect 9090 24390 9150 25230
rect 9570 25110 9630 25320
rect 9840 25290 9900 25320
rect 9780 25230 9900 25290
rect 9990 25290 10050 25320
rect 10350 25290 10410 25320
rect 9570 24480 9630 24990
rect 9780 24810 9840 25230
rect 9990 25170 10020 25290
rect 10260 25230 10410 25290
rect 10500 25290 10560 25320
rect 10770 25290 10830 25320
rect 10500 25230 10830 25290
rect 10260 25050 10320 25230
rect 10770 25110 10830 25230
rect 10080 24990 10320 25050
rect 9810 24570 9870 24690
rect 9810 24510 9900 24570
rect 9840 24480 9900 24510
rect 9990 24480 10050 24930
rect 10500 24720 10560 24990
rect 10350 24660 10560 24720
rect 10350 24480 10410 24660
rect 10770 24570 10830 24990
rect 10500 24510 10830 24570
rect 10500 24480 10560 24510
rect 10770 24480 10830 24510
rect 12210 24480 12270 25620
rect 13890 25530 13950 25620
rect 13890 25410 13980 25530
rect 12450 24990 12510 25320
rect 12600 25290 12660 25320
rect 12600 25230 12840 25290
rect 12450 24870 12540 24990
rect 12450 24480 12510 24870
rect 12780 24690 12840 25230
rect 12690 24480 12750 24630
rect 9090 24270 9180 24390
rect 9090 23880 9150 24270
rect 13890 23880 13950 25410
rect 30450 25530 30510 25620
rect 30450 25410 30540 25530
rect 15090 24210 15150 25320
rect 15330 24930 15390 25320
rect 15570 25170 15630 25320
rect 20940 25290 21000 25320
rect 20850 25230 21000 25290
rect 21090 25230 21150 25320
rect 23250 25230 23310 25320
rect 23400 25290 23460 25320
rect 25650 25290 25710 25320
rect 25920 25290 25980 25320
rect 23400 25230 23550 25290
rect 15330 24810 15420 24930
rect 15330 24570 15390 24810
rect 15660 24690 15720 25110
rect 15570 24630 15720 24690
rect 15330 24510 15480 24570
rect 15420 24480 15480 24510
rect 15570 24480 15630 24630
rect 15180 23880 15240 24150
rect 20850 24390 20910 25230
rect 20820 24270 20910 24390
rect 20850 23880 20910 24270
rect 21090 25110 21180 25230
rect 23220 25110 23310 25230
rect 21090 23880 21150 25110
rect 23250 23880 23310 25110
rect 23490 24390 23550 25230
rect 25650 25230 25980 25290
rect 26070 25290 26130 25320
rect 26430 25290 26490 25320
rect 26070 25230 26220 25290
rect 25650 25110 25710 25230
rect 26160 25050 26220 25230
rect 26460 25170 26490 25290
rect 26580 25290 26640 25320
rect 26580 25230 26700 25290
rect 26160 24990 26400 25050
rect 25650 24570 25710 24990
rect 25920 24720 25980 24990
rect 25920 24660 26130 24720
rect 25650 24510 25980 24570
rect 25650 24480 25710 24510
rect 25920 24480 25980 24510
rect 26070 24480 26130 24660
rect 26430 24480 26490 24930
rect 26640 24810 26700 25230
rect 26850 25110 26910 25320
rect 26610 24570 26670 24690
rect 26580 24510 26670 24570
rect 26580 24480 26640 24510
rect 26850 24480 26910 24990
rect 23490 24270 23580 24390
rect 23490 23880 23550 24270
rect 28050 24210 28110 25320
rect 28290 24930 28350 25320
rect 28530 25170 28590 25320
rect 28290 24810 28380 24930
rect 28290 24570 28350 24810
rect 28620 24690 28680 25110
rect 28530 24630 28680 24690
rect 28290 24510 28440 24570
rect 28380 24480 28440 24510
rect 28530 24480 28590 24630
rect 28140 23880 28200 24150
rect 30450 23880 30510 25410
rect 32370 25530 32430 25620
rect 32370 25410 32460 25530
rect 31170 24210 31230 25320
rect 31410 24930 31470 25320
rect 31650 25170 31710 25320
rect 31410 24810 31500 24930
rect 31410 24570 31470 24810
rect 31740 24690 31800 25110
rect 31650 24630 31800 24690
rect 31410 24510 31560 24570
rect 31500 24480 31560 24510
rect 31650 24480 31710 24630
rect 31260 23880 31320 24150
rect 32370 23880 32430 25410
rect 43410 25530 43470 25620
rect 43380 25410 43470 25530
rect 33330 25230 33390 25320
rect 33480 25290 33540 25320
rect 33480 25230 33630 25290
rect 34770 25230 34830 25320
rect 34920 25290 34980 25320
rect 34920 25230 35070 25290
rect 36210 25230 36270 25320
rect 36360 25290 36420 25320
rect 36360 25230 36510 25290
rect 37650 25230 37710 25320
rect 37800 25290 37860 25320
rect 37800 25230 37950 25290
rect 39090 25230 39150 25320
rect 39240 25290 39300 25320
rect 39240 25230 39390 25290
rect 40530 25230 40590 25320
rect 40680 25290 40740 25320
rect 40680 25230 40830 25290
rect 41970 25230 42030 25320
rect 42120 25290 42180 25320
rect 42120 25230 42270 25290
rect 33300 25110 33390 25230
rect 33330 23880 33390 25110
rect 33570 24390 33630 25230
rect 34740 25110 34830 25230
rect 33570 24270 33660 24390
rect 33570 23880 33630 24270
rect 34770 23880 34830 25110
rect 35010 24390 35070 25230
rect 36180 25110 36270 25230
rect 35010 24270 35100 24390
rect 35010 23880 35070 24270
rect 36210 23880 36270 25110
rect 36450 24390 36510 25230
rect 37620 25110 37710 25230
rect 36450 24270 36540 24390
rect 36450 23880 36510 24270
rect 37650 23880 37710 25110
rect 37890 24390 37950 25230
rect 39060 25110 39150 25230
rect 37890 24270 37980 24390
rect 37890 23880 37950 24270
rect 39090 23880 39150 25110
rect 39330 24390 39390 25230
rect 40500 25110 40590 25230
rect 39330 24270 39420 24390
rect 39330 23880 39390 24270
rect 40530 23880 40590 25110
rect 40770 24390 40830 25230
rect 41940 25110 42030 25230
rect 40770 24270 40860 24390
rect 40770 23880 40830 24270
rect 41970 23880 42030 25110
rect 42210 24390 42270 25230
rect 43410 24480 43470 25410
rect 43650 24690 43710 25620
rect 44610 25530 44670 25620
rect 44580 25410 44670 25530
rect 43650 24570 43740 24690
rect 43560 24510 43710 24570
rect 43560 24480 43620 24510
rect 42210 24270 42300 24390
rect 42210 23880 42270 24270
rect 44610 23880 44670 25410
rect 47970 25110 48030 25320
rect 48240 25290 48300 25320
rect 48180 25230 48300 25290
rect 48390 25290 48450 25320
rect 48750 25290 48810 25320
rect 47970 24480 48030 24990
rect 48180 24810 48240 25230
rect 48390 25170 48420 25290
rect 48660 25230 48810 25290
rect 48900 25290 48960 25320
rect 49170 25290 49230 25320
rect 48900 25230 49230 25290
rect 48660 25050 48720 25230
rect 49170 25110 49230 25230
rect 48480 24990 48720 25050
rect 48210 24570 48270 24690
rect 48210 24510 48300 24570
rect 48240 24480 48300 24510
rect 48390 24480 48450 24930
rect 48900 24720 48960 24990
rect 48750 24660 48960 24720
rect 48750 24480 48810 24660
rect 49170 24570 49230 24990
rect 48900 24510 49230 24570
rect 48900 24480 48960 24510
rect 49170 24480 49230 24510
rect 5490 23220 5550 23280
rect 5760 23220 5820 23280
rect 5910 23220 5970 23280
rect 6270 23220 6330 23280
rect 6420 23220 6480 23280
rect 6690 23220 6750 23280
rect 7170 23220 7230 23280
rect 7410 23220 7470 23280
rect 7980 23220 8040 23280
rect 8220 23220 8280 23280
rect 8370 23220 8430 23280
rect 8850 23220 8910 23280
rect 9090 23220 9150 23280
rect 9570 23220 9630 23280
rect 9840 23220 9900 23280
rect 9990 23220 10050 23280
rect 10350 23220 10410 23280
rect 10500 23220 10560 23280
rect 10770 23220 10830 23280
rect 12210 23220 12270 23280
rect 12450 23220 12510 23280
rect 12690 23220 12750 23280
rect 13890 23220 13950 23280
rect 15180 23220 15240 23280
rect 15420 23220 15480 23280
rect 15570 23220 15630 23280
rect 20850 23220 20910 23280
rect 21090 23220 21150 23280
rect 23250 23220 23310 23280
rect 23490 23220 23550 23280
rect 25650 23220 25710 23280
rect 25920 23220 25980 23280
rect 26070 23220 26130 23280
rect 26430 23220 26490 23280
rect 26580 23220 26640 23280
rect 26850 23220 26910 23280
rect 28140 23220 28200 23280
rect 28380 23220 28440 23280
rect 28530 23220 28590 23280
rect 30450 23220 30510 23280
rect 31260 23220 31320 23280
rect 31500 23220 31560 23280
rect 31650 23220 31710 23280
rect 32370 23220 32430 23280
rect 33330 23220 33390 23280
rect 33570 23220 33630 23280
rect 34770 23220 34830 23280
rect 35010 23220 35070 23280
rect 36210 23220 36270 23280
rect 36450 23220 36510 23280
rect 37650 23220 37710 23280
rect 37890 23220 37950 23280
rect 39090 23220 39150 23280
rect 39330 23220 39390 23280
rect 40530 23220 40590 23280
rect 40770 23220 40830 23280
rect 41970 23220 42030 23280
rect 42210 23220 42270 23280
rect 43410 23220 43470 23280
rect 43560 23220 43620 23280
rect 44610 23220 44670 23280
rect 47970 23220 48030 23280
rect 48240 23220 48300 23280
rect 48390 23220 48450 23280
rect 48750 23220 48810 23280
rect 48900 23220 48960 23280
rect 49170 23220 49230 23280
rect 5490 22920 5550 22980
rect 5760 22920 5820 22980
rect 5910 22920 5970 22980
rect 6270 22920 6330 22980
rect 6420 22920 6480 22980
rect 6690 22920 6750 22980
rect 8370 22920 8430 22980
rect 8610 22920 8670 22980
rect 9810 22920 9870 22980
rect 10050 22920 10110 22980
rect 11340 22920 11400 22980
rect 11580 22920 11640 22980
rect 11730 22920 11790 22980
rect 14370 22920 14430 22980
rect 14640 22920 14700 22980
rect 14790 22920 14850 22980
rect 15150 22920 15210 22980
rect 15300 22920 15360 22980
rect 15570 22920 15630 22980
rect 17010 22920 17070 22980
rect 18210 22920 18270 22980
rect 18450 22920 18510 22980
rect 18930 22920 18990 22980
rect 19200 22920 19260 22980
rect 19350 22920 19410 22980
rect 19710 22920 19770 22980
rect 19860 22920 19920 22980
rect 20130 22920 20190 22980
rect 20610 22920 20670 22980
rect 20880 22920 20940 22980
rect 21030 22920 21090 22980
rect 21390 22920 21450 22980
rect 21540 22920 21600 22980
rect 21810 22920 21870 22980
rect 22380 22920 22440 22980
rect 22620 22920 22680 22980
rect 22770 22920 22830 22980
rect 25170 22920 25230 22980
rect 26460 22920 26520 22980
rect 26700 22920 26760 22980
rect 26850 22920 26910 22980
rect 28140 22920 28200 22980
rect 28380 22920 28440 22980
rect 28530 22920 28590 22980
rect 29250 22920 29310 22980
rect 29490 22920 29550 22980
rect 30450 22920 30510 22980
rect 30600 22920 30660 22980
rect 30840 22920 30900 22980
rect 32130 22920 32190 22980
rect 32370 22920 32430 22980
rect 33330 22920 33390 22980
rect 33570 22920 33630 22980
rect 34770 22920 34830 22980
rect 35010 22920 35070 22980
rect 35970 22920 36030 22980
rect 36210 22920 36270 22980
rect 36930 22920 36990 22980
rect 37200 22920 37260 22980
rect 37350 22920 37410 22980
rect 37710 22920 37770 22980
rect 37860 22920 37920 22980
rect 38130 22920 38190 22980
rect 39180 22920 39240 22980
rect 39420 22920 39480 22980
rect 39570 22920 39630 22980
rect 40530 22920 40590 22980
rect 40770 22920 40830 22980
rect 41820 22920 41880 22980
rect 42060 22920 42120 22980
rect 42210 22920 42270 22980
rect 43410 22920 43470 22980
rect 43560 22920 43620 22980
rect 44370 22920 44430 22980
rect 44640 22920 44700 22980
rect 44790 22920 44850 22980
rect 45150 22920 45210 22980
rect 45300 22920 45360 22980
rect 45570 22920 45630 22980
rect 46050 22920 46110 22980
rect 46320 22920 46380 22980
rect 46470 22920 46530 22980
rect 46830 22920 46890 22980
rect 46980 22920 47040 22980
rect 47250 22920 47310 22980
rect 47730 22920 47790 22980
rect 48930 22920 48990 22980
rect 49170 22920 49230 22980
rect 49410 22920 49470 22980
rect 49650 22920 49710 22980
rect 5490 21210 5550 21720
rect 5760 21690 5820 21720
rect 5730 21630 5820 21690
rect 5730 21510 5790 21630
rect 5490 20880 5550 21090
rect 5700 20970 5760 21390
rect 5910 21270 5970 21720
rect 6270 21540 6330 21720
rect 6420 21690 6480 21720
rect 6690 21690 6750 21720
rect 6420 21630 6750 21690
rect 6270 21480 6480 21540
rect 6420 21210 6480 21480
rect 6690 21210 6750 21630
rect 6000 21150 6240 21210
rect 5700 20910 5820 20970
rect 5760 20880 5820 20910
rect 5910 20910 5940 21030
rect 6180 20970 6240 21150
rect 8370 21090 8430 22320
rect 6690 20970 6750 21090
rect 8340 20970 8430 21090
rect 8610 21930 8670 22320
rect 8610 21810 8700 21930
rect 8610 20970 8670 21810
rect 9810 21090 9870 22320
rect 9780 20970 9870 21090
rect 10050 21930 10110 22320
rect 11340 22050 11400 22320
rect 10050 21810 10140 21930
rect 10050 20970 10110 21810
rect 6180 20910 6330 20970
rect 5910 20880 5970 20910
rect 6270 20880 6330 20910
rect 6420 20910 6750 20970
rect 6420 20880 6480 20910
rect 6690 20880 6750 20910
rect 8370 20880 8430 20970
rect 8520 20910 8670 20970
rect 8520 20880 8580 20910
rect 9810 20880 9870 20970
rect 9960 20910 10110 20970
rect 9960 20880 10020 20910
rect 11250 20880 11310 21990
rect 11580 21690 11640 21720
rect 11490 21630 11640 21690
rect 11490 21390 11550 21630
rect 11730 21570 11790 21720
rect 11730 21510 11880 21570
rect 11490 21270 11580 21390
rect 11490 20880 11550 21270
rect 11820 21090 11880 21510
rect 14370 21210 14430 21720
rect 14640 21690 14700 21720
rect 14610 21630 14700 21690
rect 14610 21510 14670 21630
rect 11730 20880 11790 21030
rect 14370 20880 14430 21090
rect 14580 20970 14640 21390
rect 14790 21270 14850 21720
rect 15150 21540 15210 21720
rect 15300 21690 15360 21720
rect 15570 21690 15630 21720
rect 15300 21630 15630 21690
rect 15150 21480 15360 21540
rect 15300 21210 15360 21480
rect 15570 21210 15630 21630
rect 14880 21150 15120 21210
rect 14580 20910 14700 20970
rect 14640 20880 14700 20910
rect 14790 20910 14820 21030
rect 15060 20970 15120 21150
rect 15570 20970 15630 21090
rect 15060 20910 15210 20970
rect 14790 20880 14850 20910
rect 15150 20880 15210 20910
rect 15300 20910 15630 20970
rect 15300 20880 15360 20910
rect 15570 20880 15630 20910
rect 17010 20790 17070 22320
rect 18210 21090 18270 22320
rect 18180 20970 18270 21090
rect 18450 21930 18510 22320
rect 18450 21810 18540 21930
rect 18450 20970 18510 21810
rect 22380 22050 22440 22320
rect 18930 21690 18990 21720
rect 19200 21690 19260 21720
rect 18930 21630 19260 21690
rect 18930 21210 18990 21630
rect 19350 21540 19410 21720
rect 19200 21480 19410 21540
rect 19200 21210 19260 21480
rect 19710 21270 19770 21720
rect 19860 21690 19920 21720
rect 19860 21630 19950 21690
rect 19890 21510 19950 21630
rect 19440 21150 19680 21210
rect 18210 20880 18270 20970
rect 18360 20910 18510 20970
rect 18930 20970 18990 21090
rect 19440 20970 19500 21150
rect 18930 20910 19260 20970
rect 18360 20880 18420 20910
rect 18930 20880 18990 20910
rect 19200 20880 19260 20910
rect 19350 20910 19500 20970
rect 19740 20910 19770 21030
rect 19920 20970 19980 21390
rect 20130 21210 20190 21720
rect 20610 21690 20670 21720
rect 20880 21690 20940 21720
rect 20610 21630 20940 21690
rect 20610 21210 20670 21630
rect 21030 21540 21090 21720
rect 20880 21480 21090 21540
rect 20880 21210 20940 21480
rect 21390 21270 21450 21720
rect 21540 21690 21600 21720
rect 21540 21630 21630 21690
rect 21570 21510 21630 21630
rect 21120 21150 21360 21210
rect 19350 20880 19410 20910
rect 19710 20880 19770 20910
rect 19860 20910 19980 20970
rect 19860 20880 19920 20910
rect 20130 20880 20190 21090
rect 20610 20970 20670 21090
rect 21120 20970 21180 21150
rect 20610 20910 20940 20970
rect 20610 20880 20670 20910
rect 20880 20880 20940 20910
rect 21030 20910 21180 20970
rect 21420 20910 21450 21030
rect 21600 20970 21660 21390
rect 21810 21210 21870 21720
rect 21030 20880 21090 20910
rect 21390 20880 21450 20910
rect 21540 20910 21660 20970
rect 21540 20880 21600 20910
rect 21810 20880 21870 21090
rect 22290 20880 22350 21990
rect 22620 21690 22680 21720
rect 22530 21630 22680 21690
rect 22530 21390 22590 21630
rect 22770 21570 22830 21720
rect 22770 21510 22920 21570
rect 22530 21270 22620 21390
rect 22530 20880 22590 21270
rect 22860 21090 22920 21510
rect 22770 20880 22830 21030
rect 17010 20670 17100 20790
rect 17010 20580 17070 20670
rect 25170 20790 25230 22320
rect 26460 22050 26520 22320
rect 26370 20880 26430 21990
rect 28140 22050 28200 22320
rect 26700 21690 26760 21720
rect 26610 21630 26760 21690
rect 26610 21390 26670 21630
rect 26850 21570 26910 21720
rect 26850 21510 27000 21570
rect 26610 21270 26700 21390
rect 26610 20880 26670 21270
rect 26940 21090 27000 21510
rect 26850 20880 26910 21030
rect 28050 20880 28110 21990
rect 28380 21690 28440 21720
rect 28290 21630 28440 21690
rect 28290 21390 28350 21630
rect 28530 21570 28590 21720
rect 28530 21510 28680 21570
rect 28290 21270 28380 21390
rect 28290 20880 28350 21270
rect 28620 21090 28680 21510
rect 29250 21090 29310 22320
rect 28530 20880 28590 21030
rect 29220 20970 29310 21090
rect 29490 21930 29550 22320
rect 29490 21810 29580 21930
rect 29490 20970 29550 21810
rect 30840 22050 30900 22320
rect 30450 21570 30510 21720
rect 30600 21690 30660 21720
rect 30600 21630 30750 21690
rect 30360 21510 30510 21570
rect 30360 21090 30420 21510
rect 30690 21390 30750 21630
rect 30660 21270 30750 21390
rect 29250 20880 29310 20970
rect 29400 20910 29550 20970
rect 29400 20880 29460 20910
rect 30450 20880 30510 21030
rect 30690 20880 30750 21270
rect 30930 20880 30990 21990
rect 32130 21090 32190 22320
rect 32100 20970 32190 21090
rect 32370 21930 32430 22320
rect 32370 21810 32460 21930
rect 32370 20970 32430 21810
rect 33330 21090 33390 22320
rect 33300 20970 33390 21090
rect 33570 21930 33630 22320
rect 33570 21810 33660 21930
rect 33570 20970 33630 21810
rect 34770 21090 34830 22320
rect 34740 20970 34830 21090
rect 35010 21930 35070 22320
rect 35010 21810 35100 21930
rect 35010 20970 35070 21810
rect 35970 21090 36030 22320
rect 35940 20970 36030 21090
rect 36210 21930 36270 22320
rect 36210 21810 36300 21930
rect 36210 20970 36270 21810
rect 39180 22050 39240 22320
rect 36930 21210 36990 21720
rect 37200 21690 37260 21720
rect 37170 21630 37260 21690
rect 37170 21510 37230 21630
rect 32130 20880 32190 20970
rect 32280 20910 32430 20970
rect 32280 20880 32340 20910
rect 33330 20880 33390 20970
rect 33480 20910 33630 20970
rect 33480 20880 33540 20910
rect 34770 20880 34830 20970
rect 34920 20910 35070 20970
rect 34920 20880 34980 20910
rect 35970 20880 36030 20970
rect 36120 20910 36270 20970
rect 36120 20880 36180 20910
rect 36930 20880 36990 21090
rect 37140 20970 37200 21390
rect 37350 21270 37410 21720
rect 37710 21540 37770 21720
rect 37860 21690 37920 21720
rect 38130 21690 38190 21720
rect 37860 21630 38190 21690
rect 37710 21480 37920 21540
rect 37860 21210 37920 21480
rect 38130 21210 38190 21630
rect 37440 21150 37680 21210
rect 37140 20910 37260 20970
rect 37200 20880 37260 20910
rect 37350 20910 37380 21030
rect 37620 20970 37680 21150
rect 38130 20970 38190 21090
rect 37620 20910 37770 20970
rect 37350 20880 37410 20910
rect 37710 20880 37770 20910
rect 37860 20910 38190 20970
rect 37860 20880 37920 20910
rect 38130 20880 38190 20910
rect 39090 20880 39150 21990
rect 39420 21690 39480 21720
rect 39330 21630 39480 21690
rect 39330 21390 39390 21630
rect 39570 21570 39630 21720
rect 39570 21510 39720 21570
rect 39330 21270 39420 21390
rect 39330 20880 39390 21270
rect 39660 21090 39720 21510
rect 40530 21090 40590 22320
rect 39570 20880 39630 21030
rect 40500 20970 40590 21090
rect 40770 21930 40830 22320
rect 41820 22050 41880 22320
rect 40770 21810 40860 21930
rect 40770 20970 40830 21810
rect 40530 20880 40590 20970
rect 40680 20910 40830 20970
rect 40680 20880 40740 20910
rect 41730 20880 41790 21990
rect 42060 21690 42120 21720
rect 41970 21630 42120 21690
rect 41970 21390 42030 21630
rect 42210 21570 42270 21720
rect 42210 21510 42360 21570
rect 41970 21270 42060 21390
rect 41970 20880 42030 21270
rect 42300 21090 42360 21510
rect 42210 20880 42270 21030
rect 25140 20670 25230 20790
rect 25170 20580 25230 20670
rect 43410 20790 43470 21720
rect 43560 21690 43620 21720
rect 43560 21630 43710 21690
rect 43380 20670 43470 20790
rect 43410 20580 43470 20670
rect 43650 21510 43740 21630
rect 43650 20580 43710 21510
rect 44370 21210 44430 21720
rect 44640 21690 44700 21720
rect 44610 21630 44700 21690
rect 44610 21510 44670 21630
rect 44370 20880 44430 21090
rect 44580 20970 44640 21390
rect 44790 21270 44850 21720
rect 45150 21540 45210 21720
rect 45300 21690 45360 21720
rect 45570 21690 45630 21720
rect 45300 21630 45630 21690
rect 45150 21480 45360 21540
rect 45300 21210 45360 21480
rect 45570 21210 45630 21630
rect 46050 21690 46110 21720
rect 46320 21690 46380 21720
rect 46050 21630 46380 21690
rect 46050 21210 46110 21630
rect 46470 21540 46530 21720
rect 46320 21480 46530 21540
rect 46320 21210 46380 21480
rect 46830 21270 46890 21720
rect 46980 21690 47040 21720
rect 46980 21630 47070 21690
rect 47010 21510 47070 21630
rect 44880 21150 45120 21210
rect 44580 20910 44700 20970
rect 44640 20880 44700 20910
rect 44790 20910 44820 21030
rect 45060 20970 45120 21150
rect 46560 21150 46800 21210
rect 45570 20970 45630 21090
rect 45060 20910 45210 20970
rect 44790 20880 44850 20910
rect 45150 20880 45210 20910
rect 45300 20910 45630 20970
rect 45300 20880 45360 20910
rect 45570 20880 45630 20910
rect 46050 20970 46110 21090
rect 46560 20970 46620 21150
rect 46050 20910 46380 20970
rect 46050 20880 46110 20910
rect 46320 20880 46380 20910
rect 46470 20910 46620 20970
rect 46860 20910 46890 21030
rect 47040 20970 47100 21390
rect 47250 21210 47310 21720
rect 46470 20880 46530 20910
rect 46830 20880 46890 20910
rect 46980 20910 47100 20970
rect 46980 20880 47040 20910
rect 47250 20880 47310 21090
rect 47730 20790 47790 22320
rect 48930 21690 48990 21720
rect 48870 21630 48990 21690
rect 48900 21510 48930 21630
rect 48870 21030 48930 21510
rect 49170 21300 49230 21720
rect 49410 21690 49470 21720
rect 49410 21630 49500 21690
rect 49170 21270 49200 21300
rect 48870 20970 48990 21030
rect 49140 20970 49200 21270
rect 48930 20880 48990 20970
rect 49080 20910 49200 20970
rect 49080 20880 49140 20910
rect 49440 20880 49500 21630
rect 49650 21570 49710 21720
rect 49740 20970 49800 21510
rect 49590 20910 49800 20970
rect 49590 20880 49650 20910
rect 47700 20670 47790 20790
rect 47730 20580 47790 20670
rect 5490 20220 5550 20280
rect 5760 20220 5820 20280
rect 5910 20220 5970 20280
rect 6270 20220 6330 20280
rect 6420 20220 6480 20280
rect 6690 20220 6750 20280
rect 8370 20220 8430 20280
rect 8520 20220 8580 20280
rect 9810 20220 9870 20280
rect 9960 20220 10020 20280
rect 11250 20220 11310 20280
rect 11490 20220 11550 20280
rect 11730 20220 11790 20280
rect 14370 20220 14430 20280
rect 14640 20220 14700 20280
rect 14790 20220 14850 20280
rect 15150 20220 15210 20280
rect 15300 20220 15360 20280
rect 15570 20220 15630 20280
rect 17010 20220 17070 20280
rect 18210 20220 18270 20280
rect 18360 20220 18420 20280
rect 18930 20220 18990 20280
rect 19200 20220 19260 20280
rect 19350 20220 19410 20280
rect 19710 20220 19770 20280
rect 19860 20220 19920 20280
rect 20130 20220 20190 20280
rect 20610 20220 20670 20280
rect 20880 20220 20940 20280
rect 21030 20220 21090 20280
rect 21390 20220 21450 20280
rect 21540 20220 21600 20280
rect 21810 20220 21870 20280
rect 22290 20220 22350 20280
rect 22530 20220 22590 20280
rect 22770 20220 22830 20280
rect 25170 20220 25230 20280
rect 26370 20220 26430 20280
rect 26610 20220 26670 20280
rect 26850 20220 26910 20280
rect 28050 20220 28110 20280
rect 28290 20220 28350 20280
rect 28530 20220 28590 20280
rect 29250 20220 29310 20280
rect 29400 20220 29460 20280
rect 30450 20220 30510 20280
rect 30690 20220 30750 20280
rect 30930 20220 30990 20280
rect 32130 20220 32190 20280
rect 32280 20220 32340 20280
rect 33330 20220 33390 20280
rect 33480 20220 33540 20280
rect 34770 20220 34830 20280
rect 34920 20220 34980 20280
rect 35970 20220 36030 20280
rect 36120 20220 36180 20280
rect 36930 20220 36990 20280
rect 37200 20220 37260 20280
rect 37350 20220 37410 20280
rect 37710 20220 37770 20280
rect 37860 20220 37920 20280
rect 38130 20220 38190 20280
rect 39090 20220 39150 20280
rect 39330 20220 39390 20280
rect 39570 20220 39630 20280
rect 40530 20220 40590 20280
rect 40680 20220 40740 20280
rect 41730 20220 41790 20280
rect 41970 20220 42030 20280
rect 42210 20220 42270 20280
rect 43410 20220 43470 20280
rect 43650 20220 43710 20280
rect 44370 20220 44430 20280
rect 44640 20220 44700 20280
rect 44790 20220 44850 20280
rect 45150 20220 45210 20280
rect 45300 20220 45360 20280
rect 45570 20220 45630 20280
rect 46050 20220 46110 20280
rect 46320 20220 46380 20280
rect 46470 20220 46530 20280
rect 46830 20220 46890 20280
rect 46980 20220 47040 20280
rect 47250 20220 47310 20280
rect 47730 20220 47790 20280
rect 48930 20220 48990 20280
rect 49080 20220 49140 20280
rect 49440 20220 49500 20280
rect 49590 20220 49650 20280
rect 5730 19920 5790 19980
rect 5970 19920 6030 19980
rect 6210 19920 6270 19980
rect 9090 19920 9150 19980
rect 9360 19920 9420 19980
rect 9510 19920 9570 19980
rect 9870 19920 9930 19980
rect 10020 19920 10080 19980
rect 10290 19920 10350 19980
rect 11730 19920 11790 19980
rect 12000 19920 12060 19980
rect 12150 19920 12210 19980
rect 12510 19920 12570 19980
rect 12660 19920 12720 19980
rect 12930 19920 12990 19980
rect 13650 19920 13710 19980
rect 13920 19920 13980 19980
rect 14070 19920 14130 19980
rect 14430 19920 14490 19980
rect 14580 19920 14640 19980
rect 14850 19920 14910 19980
rect 15660 19920 15720 19980
rect 15810 19920 15870 19980
rect 16050 19920 16110 19980
rect 17970 19920 18030 19980
rect 18210 19920 18270 19980
rect 18450 19920 18510 19980
rect 19650 19920 19710 19980
rect 19800 19920 19860 19980
rect 21090 19920 21150 19980
rect 21240 19920 21300 19980
rect 22290 19920 22350 19980
rect 22440 19920 22500 19980
rect 23730 19920 23790 19980
rect 23880 19920 23940 19980
rect 24690 19920 24750 19980
rect 24960 19920 25020 19980
rect 25110 19920 25170 19980
rect 25470 19920 25530 19980
rect 25620 19920 25680 19980
rect 25890 19920 25950 19980
rect 26370 19920 26430 19980
rect 26610 19920 26670 19980
rect 26850 19920 26910 19980
rect 27330 19920 27390 19980
rect 28530 19920 28590 19980
rect 28770 19920 28830 19980
rect 29010 19920 29070 19980
rect 30690 19920 30750 19980
rect 30840 19920 30900 19980
rect 32130 19920 32190 19980
rect 32280 19920 32340 19980
rect 33330 19920 33390 19980
rect 33570 19920 33630 19980
rect 33810 19920 33870 19980
rect 35970 19920 36030 19980
rect 36120 19920 36180 19980
rect 36930 19920 36990 19980
rect 37170 19920 37230 19980
rect 37320 19920 37380 19980
rect 38130 19920 38190 19980
rect 38280 19920 38340 19980
rect 39090 19920 39150 19980
rect 39240 19920 39300 19980
rect 40530 19920 40590 19980
rect 40680 19920 40740 19980
rect 41730 19920 41790 19980
rect 42990 19920 43050 19980
rect 43140 19920 43200 19980
rect 43500 19920 43560 19980
rect 43650 19920 43710 19980
rect 44610 19920 44670 19980
rect 44850 19920 44910 19980
rect 45090 19920 45150 19980
rect 46290 19920 46350 19980
rect 46440 19920 46500 19980
rect 47730 19920 47790 19980
rect 47970 19920 48030 19980
rect 49170 19920 49230 19980
rect 49410 19920 49470 19980
rect 49650 19920 49710 19980
rect 5730 18210 5790 19320
rect 5970 18930 6030 19320
rect 6210 19170 6270 19320
rect 9090 19290 9150 19320
rect 9360 19290 9420 19320
rect 9090 19230 9420 19290
rect 9510 19290 9570 19320
rect 9870 19290 9930 19320
rect 9510 19230 9660 19290
rect 9090 19110 9150 19230
rect 5970 18810 6060 18930
rect 5970 18570 6030 18810
rect 6300 18690 6360 19110
rect 9600 19050 9660 19230
rect 9900 19170 9930 19290
rect 10020 19290 10080 19320
rect 10020 19230 10140 19290
rect 9600 18990 9840 19050
rect 6210 18630 6360 18690
rect 5970 18510 6120 18570
rect 6060 18480 6120 18510
rect 6210 18480 6270 18630
rect 9090 18570 9150 18990
rect 9360 18720 9420 18990
rect 9360 18660 9570 18720
rect 9090 18510 9420 18570
rect 9090 18480 9150 18510
rect 9360 18480 9420 18510
rect 9510 18480 9570 18660
rect 9870 18480 9930 18930
rect 10080 18810 10140 19230
rect 10290 19110 10350 19320
rect 11730 19110 11790 19320
rect 12000 19290 12060 19320
rect 11940 19230 12060 19290
rect 12150 19290 12210 19320
rect 12510 19290 12570 19320
rect 12150 19230 12180 19290
rect 10050 18570 10110 18690
rect 10020 18510 10110 18570
rect 10020 18480 10080 18510
rect 10290 18480 10350 18990
rect 11700 18600 11760 18990
rect 11940 18870 12000 19230
rect 12420 19230 12570 19290
rect 12660 19290 12720 19320
rect 12930 19290 12990 19320
rect 12660 19230 12990 19290
rect 12420 19050 12480 19230
rect 12930 19110 12990 19230
rect 13650 19110 13710 19320
rect 13920 19290 13980 19320
rect 13860 19230 13980 19290
rect 14070 19290 14130 19320
rect 14430 19290 14490 19320
rect 11700 18540 11790 18600
rect 11730 18480 11790 18540
rect 11940 18570 12000 18750
rect 12270 18990 12480 19050
rect 12270 18690 12330 18990
rect 12600 18900 12660 18990
rect 11940 18510 12060 18570
rect 12000 18480 12060 18510
rect 12150 18480 12210 18690
rect 12510 18840 12660 18900
rect 12510 18480 12570 18840
rect 12930 18570 12990 18990
rect 12660 18510 12990 18570
rect 12660 18480 12720 18510
rect 12930 18480 12990 18510
rect 13650 18480 13710 18990
rect 13860 18810 13920 19230
rect 14070 19170 14100 19290
rect 14340 19230 14490 19290
rect 14580 19290 14640 19320
rect 14850 19290 14910 19320
rect 15660 19290 15720 19320
rect 14580 19230 14910 19290
rect 14340 19050 14400 19230
rect 14850 19110 14910 19230
rect 15480 19230 15720 19290
rect 14160 18990 14400 19050
rect 13890 18570 13950 18690
rect 13890 18510 13980 18570
rect 13920 18480 13980 18510
rect 14070 18480 14130 18930
rect 14580 18720 14640 18990
rect 14430 18660 14640 18720
rect 14430 18480 14490 18660
rect 14850 18570 14910 18990
rect 15480 18690 15540 19230
rect 15810 18990 15870 19320
rect 15780 18870 15870 18990
rect 14580 18510 14910 18570
rect 14580 18480 14640 18510
rect 14850 18480 14910 18510
rect 15570 18480 15630 18630
rect 15810 18480 15870 18870
rect 16050 18480 16110 19620
rect 27330 19530 27390 19620
rect 27330 19410 27420 19530
rect 5820 17880 5880 18150
rect 17970 18210 18030 19320
rect 18210 18930 18270 19320
rect 18450 19170 18510 19320
rect 19650 19230 19710 19320
rect 19800 19290 19860 19320
rect 19800 19230 19950 19290
rect 21090 19230 21150 19320
rect 21240 19290 21300 19320
rect 21240 19230 21390 19290
rect 22290 19230 22350 19320
rect 22440 19290 22500 19320
rect 22440 19230 22590 19290
rect 23730 19230 23790 19320
rect 23880 19290 23940 19320
rect 23880 19230 24030 19290
rect 19620 19110 19710 19230
rect 18210 18810 18300 18930
rect 18210 18570 18270 18810
rect 18540 18690 18600 19110
rect 18450 18630 18600 18690
rect 18210 18510 18360 18570
rect 18300 18480 18360 18510
rect 18450 18480 18510 18630
rect 18060 17880 18120 18150
rect 19650 17880 19710 19110
rect 19890 18390 19950 19230
rect 21060 19110 21150 19230
rect 19890 18270 19980 18390
rect 19890 17880 19950 18270
rect 21090 17880 21150 19110
rect 21330 18390 21390 19230
rect 22260 19110 22350 19230
rect 21330 18270 21420 18390
rect 21330 17880 21390 18270
rect 22290 17880 22350 19110
rect 22530 18390 22590 19230
rect 23700 19110 23790 19230
rect 22530 18270 22620 18390
rect 22530 17880 22590 18270
rect 23730 17880 23790 19110
rect 23970 18390 24030 19230
rect 24690 19110 24750 19320
rect 24960 19290 25020 19320
rect 24900 19230 25020 19290
rect 25110 19290 25170 19320
rect 25470 19290 25530 19320
rect 24690 18480 24750 18990
rect 24900 18810 24960 19230
rect 25110 19170 25140 19290
rect 25380 19230 25530 19290
rect 25620 19290 25680 19320
rect 25890 19290 25950 19320
rect 25620 19230 25950 19290
rect 25380 19050 25440 19230
rect 25890 19110 25950 19230
rect 26370 19170 26430 19320
rect 25200 18990 25440 19050
rect 24930 18570 24990 18690
rect 24930 18510 25020 18570
rect 24960 18480 25020 18510
rect 25110 18480 25170 18930
rect 25620 18720 25680 18990
rect 25470 18660 25680 18720
rect 25470 18480 25530 18660
rect 25890 18570 25950 18990
rect 26280 18690 26340 19110
rect 26610 18930 26670 19320
rect 26580 18810 26670 18930
rect 26280 18630 26430 18690
rect 25620 18510 25950 18570
rect 25620 18480 25680 18510
rect 25890 18480 25950 18510
rect 26370 18480 26430 18630
rect 26610 18570 26670 18810
rect 26520 18510 26670 18570
rect 26520 18480 26580 18510
rect 23970 18270 24060 18390
rect 23970 17880 24030 18270
rect 26850 18210 26910 19320
rect 26760 17880 26820 18150
rect 27330 17880 27390 19410
rect 28530 18210 28590 19320
rect 28770 18930 28830 19320
rect 29010 19170 29070 19320
rect 30690 19230 30750 19320
rect 30840 19290 30900 19320
rect 30840 19230 30990 19290
rect 32130 19230 32190 19320
rect 32280 19290 32340 19320
rect 32280 19230 32430 19290
rect 30660 19110 30750 19230
rect 28770 18810 28860 18930
rect 28770 18570 28830 18810
rect 29100 18690 29160 19110
rect 29010 18630 29160 18690
rect 28770 18510 28920 18570
rect 28860 18480 28920 18510
rect 29010 18480 29070 18630
rect 28620 17880 28680 18150
rect 30690 17880 30750 19110
rect 30930 18390 30990 19230
rect 32100 19110 32190 19230
rect 30930 18270 31020 18390
rect 30930 17880 30990 18270
rect 32130 17880 32190 19110
rect 32370 18390 32430 19230
rect 33330 19170 33390 19320
rect 33240 18690 33300 19110
rect 33570 18930 33630 19320
rect 33540 18810 33630 18930
rect 33240 18630 33390 18690
rect 33330 18480 33390 18630
rect 33570 18570 33630 18810
rect 33480 18510 33630 18570
rect 33480 18480 33540 18510
rect 32370 18270 32460 18390
rect 32370 17880 32430 18270
rect 33810 18210 33870 19320
rect 35970 19230 36030 19320
rect 36120 19290 36180 19320
rect 36120 19230 36270 19290
rect 35940 19110 36030 19230
rect 33720 17880 33780 18150
rect 35970 17880 36030 19110
rect 36210 18390 36270 19230
rect 36930 18480 36990 19620
rect 41730 19530 41790 19620
rect 41700 19410 41790 19530
rect 37170 18990 37230 19320
rect 37320 19290 37380 19320
rect 37320 19230 37560 19290
rect 38130 19230 38190 19320
rect 38280 19290 38340 19320
rect 38280 19230 38430 19290
rect 39090 19230 39150 19320
rect 39240 19290 39300 19320
rect 39240 19230 39390 19290
rect 40530 19230 40590 19320
rect 40680 19290 40740 19320
rect 40680 19230 40830 19290
rect 37170 18870 37260 18990
rect 37170 18480 37230 18870
rect 37500 18690 37560 19230
rect 38100 19110 38190 19230
rect 37410 18480 37470 18630
rect 36210 18270 36300 18390
rect 36210 17880 36270 18270
rect 38130 17880 38190 19110
rect 38370 18390 38430 19230
rect 39060 19110 39150 19230
rect 38370 18270 38460 18390
rect 38370 17880 38430 18270
rect 39090 17880 39150 19110
rect 39330 18390 39390 19230
rect 40500 19110 40590 19230
rect 39330 18270 39420 18390
rect 39330 17880 39390 18270
rect 40530 17880 40590 19110
rect 40770 18390 40830 19230
rect 40770 18270 40860 18390
rect 40770 17880 40830 18270
rect 41730 17880 41790 19410
rect 47730 19530 47790 19620
rect 47700 19410 47790 19530
rect 42990 19290 43050 19320
rect 42840 19230 43050 19290
rect 42840 18690 42900 19230
rect 42930 18480 42990 18630
rect 43140 18570 43200 19320
rect 43500 19290 43560 19320
rect 43440 19230 43560 19290
rect 43650 19230 43710 19320
rect 43440 18930 43500 19230
rect 43650 19170 43770 19230
rect 44610 19170 44670 19320
rect 43440 18900 43470 18930
rect 43140 18510 43230 18570
rect 43170 18480 43230 18510
rect 43410 18480 43470 18900
rect 43710 18690 43770 19170
rect 44520 18690 44580 19110
rect 44850 18930 44910 19320
rect 44820 18810 44910 18930
rect 43710 18570 43740 18690
rect 44520 18630 44670 18690
rect 43650 18510 43770 18570
rect 43650 18480 43710 18510
rect 44610 18480 44670 18630
rect 44850 18570 44910 18810
rect 44760 18510 44910 18570
rect 44760 18480 44820 18510
rect 45090 18210 45150 19320
rect 46290 19230 46350 19320
rect 46440 19290 46500 19320
rect 46440 19230 46590 19290
rect 46260 19110 46350 19230
rect 45000 17880 45060 18150
rect 46290 17880 46350 19110
rect 46530 18390 46590 19230
rect 47730 18480 47790 19410
rect 47970 18690 48030 19620
rect 49170 19170 49230 19320
rect 49080 18690 49140 19110
rect 49410 18930 49470 19320
rect 49380 18810 49470 18930
rect 47970 18570 48060 18690
rect 49080 18630 49230 18690
rect 47880 18510 48030 18570
rect 47880 18480 47940 18510
rect 49170 18480 49230 18630
rect 49410 18570 49470 18810
rect 49320 18510 49470 18570
rect 49320 18480 49380 18510
rect 46530 18270 46620 18390
rect 46530 17880 46590 18270
rect 49650 18210 49710 19320
rect 49560 17880 49620 18150
rect 5820 17220 5880 17280
rect 6060 17220 6120 17280
rect 6210 17220 6270 17280
rect 9090 17220 9150 17280
rect 9360 17220 9420 17280
rect 9510 17220 9570 17280
rect 9870 17220 9930 17280
rect 10020 17220 10080 17280
rect 10290 17220 10350 17280
rect 11730 17220 11790 17280
rect 12000 17220 12060 17280
rect 12150 17220 12210 17280
rect 12510 17220 12570 17280
rect 12660 17220 12720 17280
rect 12930 17220 12990 17280
rect 13650 17220 13710 17280
rect 13920 17220 13980 17280
rect 14070 17220 14130 17280
rect 14430 17220 14490 17280
rect 14580 17220 14640 17280
rect 14850 17220 14910 17280
rect 15570 17220 15630 17280
rect 15810 17220 15870 17280
rect 16050 17220 16110 17280
rect 18060 17220 18120 17280
rect 18300 17220 18360 17280
rect 18450 17220 18510 17280
rect 19650 17220 19710 17280
rect 19890 17220 19950 17280
rect 21090 17220 21150 17280
rect 21330 17220 21390 17280
rect 22290 17220 22350 17280
rect 22530 17220 22590 17280
rect 23730 17220 23790 17280
rect 23970 17220 24030 17280
rect 24690 17220 24750 17280
rect 24960 17220 25020 17280
rect 25110 17220 25170 17280
rect 25470 17220 25530 17280
rect 25620 17220 25680 17280
rect 25890 17220 25950 17280
rect 26370 17220 26430 17280
rect 26520 17220 26580 17280
rect 26760 17220 26820 17280
rect 27330 17220 27390 17280
rect 28620 17220 28680 17280
rect 28860 17220 28920 17280
rect 29010 17220 29070 17280
rect 30690 17220 30750 17280
rect 30930 17220 30990 17280
rect 32130 17220 32190 17280
rect 32370 17220 32430 17280
rect 33330 17220 33390 17280
rect 33480 17220 33540 17280
rect 33720 17220 33780 17280
rect 35970 17220 36030 17280
rect 36210 17220 36270 17280
rect 36930 17220 36990 17280
rect 37170 17220 37230 17280
rect 37410 17220 37470 17280
rect 38130 17220 38190 17280
rect 38370 17220 38430 17280
rect 39090 17220 39150 17280
rect 39330 17220 39390 17280
rect 40530 17220 40590 17280
rect 40770 17220 40830 17280
rect 41730 17220 41790 17280
rect 42930 17220 42990 17280
rect 43170 17220 43230 17280
rect 43410 17220 43470 17280
rect 43650 17220 43710 17280
rect 44610 17220 44670 17280
rect 44760 17220 44820 17280
rect 45000 17220 45060 17280
rect 46290 17220 46350 17280
rect 46530 17220 46590 17280
rect 47730 17220 47790 17280
rect 47880 17220 47940 17280
rect 49170 17220 49230 17280
rect 49320 17220 49380 17280
rect 49560 17220 49620 17280
rect 6450 16920 6510 16980
rect 6690 16920 6750 16980
rect 7890 16920 7950 16980
rect 8160 16920 8220 16980
rect 8310 16920 8370 16980
rect 8670 16920 8730 16980
rect 8820 16920 8880 16980
rect 9090 16920 9150 16980
rect 9570 16920 9630 16980
rect 9840 16920 9900 16980
rect 9990 16920 10050 16980
rect 10350 16920 10410 16980
rect 10500 16920 10560 16980
rect 10770 16920 10830 16980
rect 11250 16920 11310 16980
rect 11520 16920 11580 16980
rect 11670 16920 11730 16980
rect 12030 16920 12090 16980
rect 12180 16920 12240 16980
rect 12450 16920 12510 16980
rect 13410 16920 13470 16980
rect 13680 16920 13740 16980
rect 13830 16920 13890 16980
rect 14190 16920 14250 16980
rect 14340 16920 14400 16980
rect 14610 16920 14670 16980
rect 15090 16920 15150 16980
rect 15360 16920 15420 16980
rect 15510 16920 15570 16980
rect 15870 16920 15930 16980
rect 16020 16920 16080 16980
rect 16290 16920 16350 16980
rect 16770 16920 16830 16980
rect 17010 16920 17070 16980
rect 17250 16920 17310 16980
rect 17730 16920 17790 16980
rect 18300 16920 18360 16980
rect 18540 16920 18600 16980
rect 18690 16920 18750 16980
rect 19410 16920 19470 16980
rect 19650 16920 19710 16980
rect 20850 16920 20910 16980
rect 21000 16920 21060 16980
rect 21240 16920 21300 16980
rect 22380 16920 22440 16980
rect 22620 16920 22680 16980
rect 22770 16920 22830 16980
rect 23730 16920 23790 16980
rect 23970 16920 24030 16980
rect 24930 16920 24990 16980
rect 25170 16920 25230 16980
rect 25890 16920 25950 16980
rect 26160 16920 26220 16980
rect 26310 16920 26370 16980
rect 26670 16920 26730 16980
rect 26820 16920 26880 16980
rect 27090 16920 27150 16980
rect 28050 16920 28110 16980
rect 28290 16920 28350 16980
rect 29250 16920 29310 16980
rect 29490 16920 29550 16980
rect 30450 16920 30510 16980
rect 30720 16920 30780 16980
rect 30870 16920 30930 16980
rect 31230 16920 31290 16980
rect 31380 16920 31440 16980
rect 31650 16920 31710 16980
rect 32370 16920 32430 16980
rect 32610 16920 32670 16980
rect 33330 16920 33390 16980
rect 33570 16920 33630 16980
rect 34770 16920 34830 16980
rect 35010 16920 35070 16980
rect 36210 16920 36270 16980
rect 36360 16920 36420 16980
rect 36600 16920 36660 16980
rect 37890 16920 37950 16980
rect 38130 16920 38190 16980
rect 38850 16920 38910 16980
rect 39120 16920 39180 16980
rect 39270 16920 39330 16980
rect 39630 16920 39690 16980
rect 39780 16920 39840 16980
rect 40050 16920 40110 16980
rect 41730 16920 41790 16980
rect 42000 16920 42060 16980
rect 42150 16920 42210 16980
rect 42510 16920 42570 16980
rect 42660 16920 42720 16980
rect 42930 16920 42990 16980
rect 44610 16920 44670 16980
rect 44760 16920 44820 16980
rect 45000 16920 45060 16980
rect 46290 16920 46350 16980
rect 46530 16920 46590 16980
rect 47730 16920 47790 16980
rect 47970 16920 48030 16980
rect 49170 16920 49230 16980
rect 49320 16920 49380 16980
rect 49560 16920 49620 16980
rect 6450 15090 6510 16320
rect 6420 14970 6510 15090
rect 6690 15930 6750 16320
rect 6690 15810 6780 15930
rect 6690 14970 6750 15810
rect 7890 15210 7950 15720
rect 8160 15690 8220 15720
rect 8130 15630 8220 15690
rect 8130 15510 8190 15630
rect 6450 14880 6510 14970
rect 6600 14910 6750 14970
rect 6600 14880 6660 14910
rect 7890 14880 7950 15090
rect 8100 14970 8160 15390
rect 8310 15270 8370 15720
rect 8670 15540 8730 15720
rect 8820 15690 8880 15720
rect 9090 15690 9150 15720
rect 8820 15630 9150 15690
rect 8670 15480 8880 15540
rect 8820 15210 8880 15480
rect 9090 15210 9150 15630
rect 9570 15210 9630 15720
rect 9840 15690 9900 15720
rect 9810 15630 9900 15690
rect 9810 15510 9870 15630
rect 8400 15150 8640 15210
rect 8100 14910 8220 14970
rect 8160 14880 8220 14910
rect 8310 14910 8340 15030
rect 8580 14970 8640 15150
rect 9090 14970 9150 15090
rect 8580 14910 8730 14970
rect 8310 14880 8370 14910
rect 8670 14880 8730 14910
rect 8820 14910 9150 14970
rect 8820 14880 8880 14910
rect 9090 14880 9150 14910
rect 9570 14880 9630 15090
rect 9780 14970 9840 15390
rect 9990 15270 10050 15720
rect 10350 15540 10410 15720
rect 10500 15690 10560 15720
rect 10770 15690 10830 15720
rect 10500 15630 10830 15690
rect 11250 15660 11310 15720
rect 11520 15690 11580 15720
rect 10350 15480 10560 15540
rect 10500 15210 10560 15480
rect 10770 15210 10830 15630
rect 11220 15600 11310 15660
rect 11460 15630 11580 15690
rect 11220 15210 11280 15600
rect 11460 15450 11520 15630
rect 11670 15510 11730 15720
rect 10080 15150 10320 15210
rect 9780 14910 9900 14970
rect 9840 14880 9900 14910
rect 9990 14910 10020 15030
rect 10260 14970 10320 15150
rect 10770 14970 10830 15090
rect 10260 14910 10410 14970
rect 9990 14880 10050 14910
rect 10350 14880 10410 14910
rect 10500 14910 10830 14970
rect 10500 14880 10560 14910
rect 10770 14880 10830 14910
rect 11250 14880 11310 15090
rect 11460 14970 11520 15330
rect 11790 15210 11850 15510
rect 12030 15360 12090 15720
rect 12180 15690 12240 15720
rect 12450 15690 12510 15720
rect 12180 15630 12510 15690
rect 13410 15660 13470 15720
rect 13680 15690 13740 15720
rect 12030 15300 12180 15360
rect 12120 15210 12180 15300
rect 12450 15210 12510 15630
rect 13380 15600 13470 15660
rect 13620 15630 13740 15690
rect 13380 15210 13440 15600
rect 13620 15450 13680 15630
rect 13830 15510 13890 15720
rect 11790 15150 12000 15210
rect 11460 14910 11580 14970
rect 11520 14880 11580 14910
rect 11670 14910 11700 14970
rect 11940 14970 12000 15150
rect 12450 14970 12510 15090
rect 11940 14910 12090 14970
rect 11670 14880 11730 14910
rect 12030 14880 12090 14910
rect 12180 14910 12510 14970
rect 12180 14880 12240 14910
rect 12450 14880 12510 14910
rect 13410 14880 13470 15090
rect 13620 14970 13680 15330
rect 13950 15210 14010 15510
rect 14190 15360 14250 15720
rect 14340 15690 14400 15720
rect 14610 15690 14670 15720
rect 14340 15630 14670 15690
rect 14190 15300 14340 15360
rect 14280 15210 14340 15300
rect 14610 15210 14670 15630
rect 15090 15210 15150 15720
rect 15360 15690 15420 15720
rect 15330 15630 15420 15690
rect 15330 15510 15390 15630
rect 13950 15150 14160 15210
rect 13620 14910 13740 14970
rect 13680 14880 13740 14910
rect 13830 14910 13860 14970
rect 14100 14970 14160 15150
rect 14610 14970 14670 15090
rect 14100 14910 14250 14970
rect 13830 14880 13890 14910
rect 14190 14880 14250 14910
rect 14340 14910 14670 14970
rect 14340 14880 14400 14910
rect 14610 14880 14670 14910
rect 15090 14880 15150 15090
rect 15300 14970 15360 15390
rect 15510 15270 15570 15720
rect 15870 15540 15930 15720
rect 16020 15690 16080 15720
rect 16290 15690 16350 15720
rect 16020 15630 16350 15690
rect 15870 15480 16080 15540
rect 16020 15210 16080 15480
rect 16290 15210 16350 15630
rect 16770 15570 16830 15720
rect 15600 15150 15840 15210
rect 15300 14910 15420 14970
rect 15360 14880 15420 14910
rect 15510 14910 15540 15030
rect 15780 14970 15840 15150
rect 16290 14970 16350 15090
rect 15780 14910 15930 14970
rect 15510 14880 15570 14910
rect 15870 14880 15930 14910
rect 16020 14910 16350 14970
rect 16680 14970 16740 15510
rect 17010 15330 17070 15720
rect 16980 15210 17070 15330
rect 16680 14910 16920 14970
rect 16020 14880 16080 14910
rect 16290 14880 16350 14910
rect 16860 14880 16920 14910
rect 17010 14880 17070 15210
rect 17250 14580 17310 15720
rect 17730 14790 17790 16320
rect 18300 16050 18360 16320
rect 18210 14880 18270 15990
rect 18540 15690 18600 15720
rect 18450 15630 18600 15690
rect 18450 15390 18510 15630
rect 18690 15570 18750 15720
rect 18690 15510 18840 15570
rect 18450 15270 18540 15390
rect 18450 14880 18510 15270
rect 18780 15090 18840 15510
rect 19410 15090 19470 16320
rect 18690 14880 18750 15030
rect 19380 14970 19470 15090
rect 19650 15930 19710 16320
rect 19650 15810 19740 15930
rect 19650 14970 19710 15810
rect 21240 16050 21300 16320
rect 22380 16050 22440 16320
rect 20850 15570 20910 15720
rect 21000 15690 21060 15720
rect 21000 15630 21150 15690
rect 20760 15510 20910 15570
rect 20760 15090 20820 15510
rect 21090 15390 21150 15630
rect 21060 15270 21150 15390
rect 19410 14880 19470 14970
rect 19560 14910 19710 14970
rect 19560 14880 19620 14910
rect 20850 14880 20910 15030
rect 21090 14880 21150 15270
rect 21330 14880 21390 15990
rect 22290 14880 22350 15990
rect 22620 15690 22680 15720
rect 22530 15630 22680 15690
rect 22530 15390 22590 15630
rect 22770 15570 22830 15720
rect 22770 15510 22920 15570
rect 22530 15270 22620 15390
rect 22530 14880 22590 15270
rect 22860 15090 22920 15510
rect 23730 15090 23790 16320
rect 22770 14880 22830 15030
rect 23700 14970 23790 15090
rect 23970 15930 24030 16320
rect 24930 15930 24990 16320
rect 23970 15810 24060 15930
rect 24900 15810 24990 15930
rect 23970 14970 24030 15810
rect 23730 14880 23790 14970
rect 23880 14910 24030 14970
rect 24930 14970 24990 15810
rect 25170 15090 25230 16320
rect 25890 15690 25950 15720
rect 26160 15690 26220 15720
rect 25890 15630 26220 15690
rect 25890 15210 25950 15630
rect 26310 15540 26370 15720
rect 26160 15480 26370 15540
rect 26160 15210 26220 15480
rect 26670 15270 26730 15720
rect 26820 15690 26880 15720
rect 26820 15630 26910 15690
rect 26850 15510 26910 15630
rect 26400 15150 26640 15210
rect 25170 14970 25260 15090
rect 25890 14970 25950 15090
rect 26400 14970 26460 15150
rect 24930 14910 25080 14970
rect 23880 14880 23940 14910
rect 25020 14880 25080 14910
rect 25170 14880 25230 14970
rect 25890 14910 26220 14970
rect 25890 14880 25950 14910
rect 26160 14880 26220 14910
rect 26310 14910 26460 14970
rect 26700 14910 26730 15030
rect 26880 14970 26940 15390
rect 27090 15210 27150 15720
rect 28050 15090 28110 16320
rect 26310 14880 26370 14910
rect 26670 14880 26730 14910
rect 26820 14910 26940 14970
rect 26820 14880 26880 14910
rect 27090 14880 27150 15090
rect 28020 14970 28110 15090
rect 28290 15930 28350 16320
rect 28290 15810 28380 15930
rect 28290 14970 28350 15810
rect 29250 15090 29310 16320
rect 29220 14970 29310 15090
rect 29490 15930 29550 16320
rect 29490 15810 29580 15930
rect 29490 14970 29550 15810
rect 32370 15930 32430 16320
rect 32340 15810 32430 15930
rect 30450 15690 30510 15720
rect 30720 15690 30780 15720
rect 30450 15630 30780 15690
rect 30450 15210 30510 15630
rect 30870 15540 30930 15720
rect 30720 15480 30930 15540
rect 30720 15210 30780 15480
rect 31230 15270 31290 15720
rect 31380 15690 31440 15720
rect 31380 15630 31470 15690
rect 31410 15510 31470 15630
rect 30960 15150 31200 15210
rect 28050 14880 28110 14970
rect 28200 14910 28350 14970
rect 28200 14880 28260 14910
rect 29250 14880 29310 14970
rect 29400 14910 29550 14970
rect 30450 14970 30510 15090
rect 30960 14970 31020 15150
rect 30450 14910 30780 14970
rect 29400 14880 29460 14910
rect 30450 14880 30510 14910
rect 30720 14880 30780 14910
rect 30870 14910 31020 14970
rect 31260 14910 31290 15030
rect 31440 14970 31500 15390
rect 31650 15210 31710 15720
rect 30870 14880 30930 14910
rect 31230 14880 31290 14910
rect 31380 14910 31500 14970
rect 31380 14880 31440 14910
rect 31650 14880 31710 15090
rect 32370 14970 32430 15810
rect 32610 15090 32670 16320
rect 33330 15090 33390 16320
rect 32610 14970 32700 15090
rect 33300 14970 33390 15090
rect 33570 15930 33630 16320
rect 33570 15810 33660 15930
rect 33570 14970 33630 15810
rect 34770 15090 34830 16320
rect 34740 14970 34830 15090
rect 35010 15930 35070 16320
rect 35010 15810 35100 15930
rect 35010 14970 35070 15810
rect 36600 16050 36660 16320
rect 36210 15570 36270 15720
rect 36360 15690 36420 15720
rect 36360 15630 36510 15690
rect 36120 15510 36270 15570
rect 36120 15090 36180 15510
rect 36450 15390 36510 15630
rect 36420 15270 36510 15390
rect 32370 14910 32520 14970
rect 32460 14880 32520 14910
rect 32610 14880 32670 14970
rect 33330 14880 33390 14970
rect 33480 14910 33630 14970
rect 33480 14880 33540 14910
rect 34770 14880 34830 14970
rect 34920 14910 35070 14970
rect 34920 14880 34980 14910
rect 36210 14880 36270 15030
rect 36450 14880 36510 15270
rect 36690 14880 36750 15990
rect 37890 15090 37950 16320
rect 37860 14970 37950 15090
rect 38130 15930 38190 16320
rect 38130 15810 38220 15930
rect 38130 14970 38190 15810
rect 45000 16050 45060 16320
rect 38850 15690 38910 15720
rect 39120 15690 39180 15720
rect 38850 15630 39180 15690
rect 38850 15210 38910 15630
rect 39270 15540 39330 15720
rect 39120 15480 39330 15540
rect 39120 15210 39180 15480
rect 39630 15270 39690 15720
rect 39780 15690 39840 15720
rect 39780 15630 39870 15690
rect 39810 15510 39870 15630
rect 39360 15150 39600 15210
rect 37890 14880 37950 14970
rect 38040 14910 38190 14970
rect 38850 14970 38910 15090
rect 39360 14970 39420 15150
rect 38850 14910 39180 14970
rect 38040 14880 38100 14910
rect 38850 14880 38910 14910
rect 39120 14880 39180 14910
rect 39270 14910 39420 14970
rect 39660 14910 39690 15030
rect 39840 14970 39900 15390
rect 40050 15210 40110 15720
rect 41730 15210 41790 15720
rect 42000 15690 42060 15720
rect 41970 15630 42060 15690
rect 41970 15510 42030 15630
rect 39270 14880 39330 14910
rect 39630 14880 39690 14910
rect 39780 14910 39900 14970
rect 39780 14880 39840 14910
rect 40050 14880 40110 15090
rect 41730 14880 41790 15090
rect 41940 14970 42000 15390
rect 42150 15270 42210 15720
rect 42510 15540 42570 15720
rect 42660 15690 42720 15720
rect 42930 15690 42990 15720
rect 42660 15630 42990 15690
rect 42510 15480 42720 15540
rect 42660 15210 42720 15480
rect 42930 15210 42990 15630
rect 44610 15570 44670 15720
rect 44760 15690 44820 15720
rect 44760 15630 44910 15690
rect 44520 15510 44670 15570
rect 42240 15150 42480 15210
rect 41940 14910 42060 14970
rect 42000 14880 42060 14910
rect 42150 14910 42180 15030
rect 42420 14970 42480 15150
rect 44520 15090 44580 15510
rect 44850 15390 44910 15630
rect 44820 15270 44910 15390
rect 42930 14970 42990 15090
rect 42420 14910 42570 14970
rect 42150 14880 42210 14910
rect 42510 14880 42570 14910
rect 42660 14910 42990 14970
rect 42660 14880 42720 14910
rect 42930 14880 42990 14910
rect 44610 14880 44670 15030
rect 44850 14880 44910 15270
rect 45090 14880 45150 15990
rect 46290 15090 46350 16320
rect 46260 14970 46350 15090
rect 46530 15930 46590 16320
rect 47730 15930 47790 16320
rect 46530 15810 46620 15930
rect 47700 15810 47790 15930
rect 46530 14970 46590 15810
rect 46290 14880 46350 14970
rect 46440 14910 46590 14970
rect 47730 14970 47790 15810
rect 47970 15090 48030 16320
rect 49560 16050 49620 16320
rect 49170 15570 49230 15720
rect 49320 15690 49380 15720
rect 49320 15630 49470 15690
rect 49080 15510 49230 15570
rect 49080 15090 49140 15510
rect 49410 15390 49470 15630
rect 49380 15270 49470 15390
rect 47970 14970 48060 15090
rect 47730 14910 47880 14970
rect 46440 14880 46500 14910
rect 47820 14880 47880 14910
rect 47970 14880 48030 14970
rect 49170 14880 49230 15030
rect 49410 14880 49470 15270
rect 49650 14880 49710 15990
rect 17730 14670 17820 14790
rect 17730 14580 17790 14670
rect 6450 14220 6510 14280
rect 6600 14220 6660 14280
rect 7890 14220 7950 14280
rect 8160 14220 8220 14280
rect 8310 14220 8370 14280
rect 8670 14220 8730 14280
rect 8820 14220 8880 14280
rect 9090 14220 9150 14280
rect 9570 14220 9630 14280
rect 9840 14220 9900 14280
rect 9990 14220 10050 14280
rect 10350 14220 10410 14280
rect 10500 14220 10560 14280
rect 10770 14220 10830 14280
rect 11250 14220 11310 14280
rect 11520 14220 11580 14280
rect 11670 14220 11730 14280
rect 12030 14220 12090 14280
rect 12180 14220 12240 14280
rect 12450 14220 12510 14280
rect 13410 14220 13470 14280
rect 13680 14220 13740 14280
rect 13830 14220 13890 14280
rect 14190 14220 14250 14280
rect 14340 14220 14400 14280
rect 14610 14220 14670 14280
rect 15090 14220 15150 14280
rect 15360 14220 15420 14280
rect 15510 14220 15570 14280
rect 15870 14220 15930 14280
rect 16020 14220 16080 14280
rect 16290 14220 16350 14280
rect 16860 14220 16920 14280
rect 17010 14220 17070 14280
rect 17250 14220 17310 14280
rect 17730 14220 17790 14280
rect 18210 14220 18270 14280
rect 18450 14220 18510 14280
rect 18690 14220 18750 14280
rect 19410 14220 19470 14280
rect 19560 14220 19620 14280
rect 20850 14220 20910 14280
rect 21090 14220 21150 14280
rect 21330 14220 21390 14280
rect 22290 14220 22350 14280
rect 22530 14220 22590 14280
rect 22770 14220 22830 14280
rect 23730 14220 23790 14280
rect 23880 14220 23940 14280
rect 25020 14220 25080 14280
rect 25170 14220 25230 14280
rect 25890 14220 25950 14280
rect 26160 14220 26220 14280
rect 26310 14220 26370 14280
rect 26670 14220 26730 14280
rect 26820 14220 26880 14280
rect 27090 14220 27150 14280
rect 28050 14220 28110 14280
rect 28200 14220 28260 14280
rect 29250 14220 29310 14280
rect 29400 14220 29460 14280
rect 30450 14220 30510 14280
rect 30720 14220 30780 14280
rect 30870 14220 30930 14280
rect 31230 14220 31290 14280
rect 31380 14220 31440 14280
rect 31650 14220 31710 14280
rect 32460 14220 32520 14280
rect 32610 14220 32670 14280
rect 33330 14220 33390 14280
rect 33480 14220 33540 14280
rect 34770 14220 34830 14280
rect 34920 14220 34980 14280
rect 36210 14220 36270 14280
rect 36450 14220 36510 14280
rect 36690 14220 36750 14280
rect 37890 14220 37950 14280
rect 38040 14220 38100 14280
rect 38850 14220 38910 14280
rect 39120 14220 39180 14280
rect 39270 14220 39330 14280
rect 39630 14220 39690 14280
rect 39780 14220 39840 14280
rect 40050 14220 40110 14280
rect 41730 14220 41790 14280
rect 42000 14220 42060 14280
rect 42150 14220 42210 14280
rect 42510 14220 42570 14280
rect 42660 14220 42720 14280
rect 42930 14220 42990 14280
rect 44610 14220 44670 14280
rect 44850 14220 44910 14280
rect 45090 14220 45150 14280
rect 46290 14220 46350 14280
rect 46440 14220 46500 14280
rect 47820 14220 47880 14280
rect 47970 14220 48030 14280
rect 49170 14220 49230 14280
rect 49410 14220 49470 14280
rect 49650 14220 49710 14280
rect 7020 13920 7080 13980
rect 7170 13920 7230 13980
rect 9090 13920 9150 13980
rect 9330 13920 9390 13980
rect 9570 13920 9630 13980
rect 9810 13920 9870 13980
rect 11010 13920 11070 13980
rect 11160 13920 11220 13980
rect 12210 13920 12270 13980
rect 12450 13920 12510 13980
rect 12690 13920 12750 13980
rect 16050 13920 16110 13980
rect 16200 13920 16260 13980
rect 16770 13920 16830 13980
rect 17010 13920 17070 13980
rect 17250 13920 17310 13980
rect 17730 13920 17790 13980
rect 18000 13920 18060 13980
rect 18150 13920 18210 13980
rect 18510 13920 18570 13980
rect 18660 13920 18720 13980
rect 18930 13920 18990 13980
rect 19410 13920 19470 13980
rect 19680 13920 19740 13980
rect 19830 13920 19890 13980
rect 20190 13920 20250 13980
rect 20340 13920 20400 13980
rect 20610 13920 20670 13980
rect 22050 13920 22110 13980
rect 22320 13920 22380 13980
rect 22470 13920 22530 13980
rect 22830 13920 22890 13980
rect 22980 13920 23040 13980
rect 23250 13920 23310 13980
rect 25170 13920 25230 13980
rect 25410 13920 25470 13980
rect 25650 13920 25710 13980
rect 26850 13920 26910 13980
rect 27000 13920 27060 13980
rect 29250 13920 29310 13980
rect 29490 13920 29550 13980
rect 29730 13920 29790 13980
rect 30450 13920 30510 13980
rect 30690 13920 30750 13980
rect 30930 13920 30990 13980
rect 32220 13920 32280 13980
rect 32370 13920 32430 13980
rect 33090 13920 33150 13980
rect 33360 13920 33420 13980
rect 33510 13920 33570 13980
rect 33870 13920 33930 13980
rect 34020 13920 34080 13980
rect 34290 13920 34350 13980
rect 34770 13920 34830 13980
rect 35010 13920 35070 13980
rect 35250 13920 35310 13980
rect 36210 13920 36270 13980
rect 36360 13920 36420 13980
rect 37650 13920 37710 13980
rect 37800 13920 37860 13980
rect 39090 13920 39150 13980
rect 39240 13920 39300 13980
rect 40290 13920 40350 13980
rect 40530 13920 40590 13980
rect 40770 13920 40830 13980
rect 41730 13920 41790 13980
rect 41880 13920 41940 13980
rect 42120 13920 42180 13980
rect 43410 13920 43470 13980
rect 43560 13920 43620 13980
rect 44610 13920 44670 13980
rect 44850 13920 44910 13980
rect 45090 13920 45150 13980
rect 46290 13920 46350 13980
rect 46440 13920 46500 13980
rect 47730 13920 47790 13980
rect 47970 13920 48030 13980
rect 48210 13920 48270 13980
rect 49500 13920 49560 13980
rect 49650 13920 49710 13980
rect 7020 13290 7080 13320
rect 6930 13230 7080 13290
rect 7170 13230 7230 13320
rect 6930 12390 6990 13230
rect 6900 12270 6990 12390
rect 6930 11880 6990 12270
rect 7170 13110 7260 13230
rect 9090 13170 9150 13320
rect 7170 11880 7230 13110
rect 9000 12690 9060 13110
rect 9330 12930 9390 13320
rect 9570 13230 9630 13320
rect 9810 13260 9870 13320
rect 9570 13170 9690 13230
rect 9810 13200 9990 13260
rect 11010 13230 11070 13320
rect 11160 13290 11220 13320
rect 11160 13230 11310 13290
rect 9300 12810 9390 12930
rect 9000 12630 9150 12690
rect 9090 12480 9150 12630
rect 9330 12570 9390 12810
rect 9240 12510 9390 12570
rect 9630 12930 9690 13170
rect 9930 12990 9990 13200
rect 10980 13110 11070 13230
rect 9630 12810 9660 12930
rect 9630 12570 9690 12810
rect 9930 12570 9990 12870
rect 9630 12510 9720 12570
rect 9240 12480 9300 12510
rect 9660 12480 9720 12510
rect 9810 12510 9990 12570
rect 9810 12480 9870 12510
rect 11010 11880 11070 13110
rect 11250 12390 11310 13230
rect 11250 12270 11340 12390
rect 11250 11880 11310 12270
rect 12210 12210 12270 13320
rect 12450 12930 12510 13320
rect 12690 13170 12750 13320
rect 16050 13230 16110 13320
rect 16200 13290 16260 13320
rect 16200 13230 16350 13290
rect 16020 13110 16110 13230
rect 12450 12810 12540 12930
rect 12450 12570 12510 12810
rect 12780 12690 12840 13110
rect 12690 12630 12840 12690
rect 12450 12510 12600 12570
rect 12540 12480 12600 12510
rect 12690 12480 12750 12630
rect 12300 11880 12360 12150
rect 16050 11880 16110 13110
rect 16290 12390 16350 13230
rect 16290 12270 16380 12390
rect 16290 11880 16350 12270
rect 16770 12210 16830 13320
rect 17010 12930 17070 13320
rect 17250 13170 17310 13320
rect 17730 13110 17790 13320
rect 18000 13290 18060 13320
rect 17940 13230 18060 13290
rect 18150 13290 18210 13320
rect 18510 13290 18570 13320
rect 17010 12810 17100 12930
rect 17010 12570 17070 12810
rect 17340 12690 17400 13110
rect 17250 12630 17400 12690
rect 17010 12510 17160 12570
rect 17100 12480 17160 12510
rect 17250 12480 17310 12630
rect 17730 12480 17790 12990
rect 17940 12810 18000 13230
rect 18150 13170 18180 13290
rect 18420 13230 18570 13290
rect 18660 13290 18720 13320
rect 18930 13290 18990 13320
rect 18660 13230 18990 13290
rect 18420 13050 18480 13230
rect 18930 13110 18990 13230
rect 19410 13290 19470 13320
rect 19680 13290 19740 13320
rect 19410 13230 19740 13290
rect 19830 13290 19890 13320
rect 20190 13290 20250 13320
rect 19830 13230 19980 13290
rect 19410 13110 19470 13230
rect 18240 12990 18480 13050
rect 19920 13050 19980 13230
rect 20220 13230 20250 13290
rect 20340 13290 20400 13320
rect 20340 13230 20460 13290
rect 19920 12990 20130 13050
rect 17970 12570 18030 12690
rect 17970 12510 18060 12570
rect 18000 12480 18060 12510
rect 18150 12480 18210 12930
rect 18660 12720 18720 12990
rect 18510 12660 18720 12720
rect 18510 12480 18570 12660
rect 18930 12570 18990 12990
rect 18660 12510 18990 12570
rect 18660 12480 18720 12510
rect 18930 12480 18990 12510
rect 19410 12570 19470 12990
rect 19740 12900 19800 12990
rect 19740 12840 19890 12900
rect 19410 12510 19740 12570
rect 19410 12480 19470 12510
rect 19680 12480 19740 12510
rect 19830 12480 19890 12840
rect 20070 12690 20130 12990
rect 20400 12870 20460 13230
rect 20610 13110 20670 13320
rect 22050 13110 22110 13320
rect 22320 13290 22380 13320
rect 22260 13230 22380 13290
rect 22470 13290 22530 13320
rect 22830 13290 22890 13320
rect 22470 13230 22500 13290
rect 20190 12480 20250 12690
rect 20400 12570 20460 12750
rect 20640 12600 20700 12990
rect 20340 12510 20460 12570
rect 20610 12540 20700 12600
rect 22020 12600 22080 12990
rect 22260 12870 22320 13230
rect 22740 13230 22890 13290
rect 22980 13290 23040 13320
rect 23250 13290 23310 13320
rect 22980 13230 23310 13290
rect 22740 13050 22800 13230
rect 23250 13110 23310 13230
rect 25170 13170 25230 13320
rect 22020 12540 22110 12600
rect 20340 12480 20400 12510
rect 20610 12480 20670 12540
rect 22050 12480 22110 12540
rect 22260 12570 22320 12750
rect 22590 12990 22800 13050
rect 22590 12690 22650 12990
rect 22920 12900 22980 12990
rect 22260 12510 22380 12570
rect 22320 12480 22380 12510
rect 22470 12480 22530 12690
rect 22830 12840 22980 12900
rect 22830 12480 22890 12840
rect 23250 12570 23310 12990
rect 25080 12690 25140 13110
rect 25410 12930 25470 13320
rect 25380 12810 25470 12930
rect 25080 12630 25230 12690
rect 22980 12510 23310 12570
rect 22980 12480 23040 12510
rect 23250 12480 23310 12510
rect 25170 12480 25230 12630
rect 25410 12570 25470 12810
rect 25320 12510 25470 12570
rect 25320 12480 25380 12510
rect 16860 11880 16920 12150
rect 25650 12210 25710 13320
rect 26850 13230 26910 13320
rect 27000 13290 27060 13320
rect 27000 13230 27150 13290
rect 26820 13110 26910 13230
rect 25560 11880 25620 12150
rect 26850 11880 26910 13110
rect 27090 12390 27150 13230
rect 29250 13170 29310 13320
rect 29160 12690 29220 13110
rect 29490 12930 29550 13320
rect 29460 12810 29550 12930
rect 29160 12630 29310 12690
rect 29250 12480 29310 12630
rect 29490 12570 29550 12810
rect 29400 12510 29550 12570
rect 29400 12480 29460 12510
rect 27090 12270 27180 12390
rect 27090 11880 27150 12270
rect 29730 12210 29790 13320
rect 30450 12210 30510 13320
rect 30690 12930 30750 13320
rect 30930 13170 30990 13320
rect 32220 13290 32280 13320
rect 32130 13230 32280 13290
rect 32370 13230 32430 13320
rect 30690 12810 30780 12930
rect 30690 12570 30750 12810
rect 31020 12690 31080 13110
rect 30930 12630 31080 12690
rect 30690 12510 30840 12570
rect 30780 12480 30840 12510
rect 30930 12480 30990 12630
rect 29640 11880 29700 12150
rect 30540 11880 30600 12150
rect 32130 12390 32190 13230
rect 32100 12270 32190 12390
rect 32130 11880 32190 12270
rect 32370 13110 32460 13230
rect 33090 13110 33150 13320
rect 33360 13290 33420 13320
rect 33300 13230 33420 13290
rect 33510 13290 33570 13320
rect 33870 13290 33930 13320
rect 32370 11880 32430 13110
rect 33090 12480 33150 12990
rect 33300 12810 33360 13230
rect 33510 13170 33540 13290
rect 33780 13230 33930 13290
rect 34020 13290 34080 13320
rect 34290 13290 34350 13320
rect 34020 13230 34350 13290
rect 33780 13050 33840 13230
rect 34290 13110 34350 13230
rect 34770 13170 34830 13320
rect 33600 12990 33840 13050
rect 33330 12570 33390 12690
rect 33330 12510 33420 12570
rect 33360 12480 33420 12510
rect 33510 12480 33570 12930
rect 34020 12720 34080 12990
rect 33870 12660 34080 12720
rect 33870 12480 33930 12660
rect 34290 12570 34350 12990
rect 34680 12690 34740 13110
rect 35010 12930 35070 13320
rect 34980 12810 35070 12930
rect 34680 12630 34830 12690
rect 34020 12510 34350 12570
rect 34020 12480 34080 12510
rect 34290 12480 34350 12510
rect 34770 12480 34830 12630
rect 35010 12570 35070 12810
rect 34920 12510 35070 12570
rect 34920 12480 34980 12510
rect 35250 12210 35310 13320
rect 36210 13230 36270 13320
rect 36360 13290 36420 13320
rect 36360 13230 36510 13290
rect 37650 13230 37710 13320
rect 37800 13290 37860 13320
rect 37800 13230 37950 13290
rect 39090 13230 39150 13320
rect 39240 13290 39300 13320
rect 39240 13230 39390 13290
rect 36180 13110 36270 13230
rect 35160 11880 35220 12150
rect 36210 11880 36270 13110
rect 36450 12390 36510 13230
rect 37620 13110 37710 13230
rect 36450 12270 36540 12390
rect 36450 11880 36510 12270
rect 37650 11880 37710 13110
rect 37890 12390 37950 13230
rect 39060 13110 39150 13230
rect 37890 12270 37980 12390
rect 37890 11880 37950 12270
rect 39090 11880 39150 13110
rect 39330 12390 39390 13230
rect 39330 12270 39420 12390
rect 39330 11880 39390 12270
rect 40290 12210 40350 13320
rect 40530 12930 40590 13320
rect 40770 13170 40830 13320
rect 40530 12810 40620 12930
rect 40530 12570 40590 12810
rect 40860 12690 40920 13110
rect 41730 12990 41790 13320
rect 41700 12870 41790 12990
rect 41880 12990 41940 13320
rect 42120 13230 42180 13620
rect 43410 13230 43470 13320
rect 43560 13290 43620 13320
rect 43560 13230 43710 13290
rect 42240 13110 42270 13200
rect 43380 13110 43470 13230
rect 41880 12930 42030 12990
rect 40770 12630 40920 12690
rect 40530 12510 40680 12570
rect 40620 12480 40680 12510
rect 40770 12480 40830 12630
rect 40380 11880 40440 12150
rect 41730 11880 41790 12870
rect 41970 12630 42030 12930
rect 41970 11880 42030 12510
rect 42210 11880 42270 13110
rect 43410 11880 43470 13110
rect 43650 12390 43710 13230
rect 44610 13170 44670 13320
rect 44520 12690 44580 13110
rect 44850 12930 44910 13320
rect 44820 12810 44910 12930
rect 44520 12630 44670 12690
rect 44610 12480 44670 12630
rect 44850 12570 44910 12810
rect 44760 12510 44910 12570
rect 44760 12480 44820 12510
rect 43650 12270 43740 12390
rect 43650 11880 43710 12270
rect 45090 12210 45150 13320
rect 46290 13230 46350 13320
rect 46440 13290 46500 13320
rect 46440 13230 46590 13290
rect 46260 13110 46350 13230
rect 45000 11880 45060 12150
rect 46290 11880 46350 13110
rect 46530 12390 46590 13230
rect 47730 13170 47790 13320
rect 47640 12690 47700 13110
rect 47970 12930 48030 13320
rect 47940 12810 48030 12930
rect 47640 12630 47790 12690
rect 47730 12480 47790 12630
rect 47970 12570 48030 12810
rect 47880 12510 48030 12570
rect 47880 12480 47940 12510
rect 46530 12270 46620 12390
rect 46530 11880 46590 12270
rect 48210 12210 48270 13320
rect 49500 13290 49560 13320
rect 49410 13230 49560 13290
rect 49650 13230 49710 13320
rect 49410 12390 49470 13230
rect 49380 12270 49470 12390
rect 48120 11880 48180 12150
rect 49410 11880 49470 12270
rect 49650 13110 49740 13230
rect 49650 11880 49710 13110
rect 6930 11220 6990 11280
rect 7170 11220 7230 11280
rect 9090 11220 9150 11280
rect 9240 11220 9300 11280
rect 9660 11220 9720 11280
rect 9810 11220 9870 11280
rect 11010 11220 11070 11280
rect 11250 11220 11310 11280
rect 12300 11220 12360 11280
rect 12540 11220 12600 11280
rect 12690 11220 12750 11280
rect 16050 11220 16110 11280
rect 16290 11220 16350 11280
rect 16860 11220 16920 11280
rect 17100 11220 17160 11280
rect 17250 11220 17310 11280
rect 17730 11220 17790 11280
rect 18000 11220 18060 11280
rect 18150 11220 18210 11280
rect 18510 11220 18570 11280
rect 18660 11220 18720 11280
rect 18930 11220 18990 11280
rect 19410 11220 19470 11280
rect 19680 11220 19740 11280
rect 19830 11220 19890 11280
rect 20190 11220 20250 11280
rect 20340 11220 20400 11280
rect 20610 11220 20670 11280
rect 22050 11220 22110 11280
rect 22320 11220 22380 11280
rect 22470 11220 22530 11280
rect 22830 11220 22890 11280
rect 22980 11220 23040 11280
rect 23250 11220 23310 11280
rect 25170 11220 25230 11280
rect 25320 11220 25380 11280
rect 25560 11220 25620 11280
rect 26850 11220 26910 11280
rect 27090 11220 27150 11280
rect 29250 11220 29310 11280
rect 29400 11220 29460 11280
rect 29640 11220 29700 11280
rect 30540 11220 30600 11280
rect 30780 11220 30840 11280
rect 30930 11220 30990 11280
rect 32130 11220 32190 11280
rect 32370 11220 32430 11280
rect 33090 11220 33150 11280
rect 33360 11220 33420 11280
rect 33510 11220 33570 11280
rect 33870 11220 33930 11280
rect 34020 11220 34080 11280
rect 34290 11220 34350 11280
rect 34770 11220 34830 11280
rect 34920 11220 34980 11280
rect 35160 11220 35220 11280
rect 36210 11220 36270 11280
rect 36450 11220 36510 11280
rect 37650 11220 37710 11280
rect 37890 11220 37950 11280
rect 39090 11220 39150 11280
rect 39330 11220 39390 11280
rect 40380 11220 40440 11280
rect 40620 11220 40680 11280
rect 40770 11220 40830 11280
rect 41730 11220 41790 11280
rect 41970 11220 42030 11280
rect 42210 11220 42270 11280
rect 43410 11220 43470 11280
rect 43650 11220 43710 11280
rect 44610 11220 44670 11280
rect 44760 11220 44820 11280
rect 45000 11220 45060 11280
rect 46290 11220 46350 11280
rect 46530 11220 46590 11280
rect 47730 11220 47790 11280
rect 47880 11220 47940 11280
rect 48120 11220 48180 11280
rect 49410 11220 49470 11280
rect 49650 11220 49710 11280
rect 5820 10920 5880 10980
rect 6060 10920 6120 10980
rect 6210 10920 6270 10980
rect 6930 10920 6990 10980
rect 7170 10920 7230 10980
rect 7890 10920 7950 10980
rect 8160 10920 8220 10980
rect 8310 10920 8370 10980
rect 8670 10920 8730 10980
rect 8820 10920 8880 10980
rect 9090 10920 9150 10980
rect 9810 10920 9870 10980
rect 10050 10920 10110 10980
rect 10290 10920 10350 10980
rect 11490 10920 11550 10980
rect 11730 10920 11790 10980
rect 13890 10920 13950 10980
rect 14160 10920 14220 10980
rect 14310 10920 14370 10980
rect 14670 10920 14730 10980
rect 14820 10920 14880 10980
rect 15090 10920 15150 10980
rect 16530 10920 16590 10980
rect 16770 10920 16830 10980
rect 17490 10920 17550 10980
rect 17760 10920 17820 10980
rect 17910 10920 17970 10980
rect 18270 10920 18330 10980
rect 18420 10920 18480 10980
rect 18690 10920 18750 10980
rect 19410 10920 19470 10980
rect 19680 10920 19740 10980
rect 19830 10920 19890 10980
rect 20190 10920 20250 10980
rect 20340 10920 20400 10980
rect 20610 10920 20670 10980
rect 21330 10920 21390 10980
rect 21570 10920 21630 10980
rect 22050 10920 22110 10980
rect 22320 10920 22380 10980
rect 22470 10920 22530 10980
rect 22830 10920 22890 10980
rect 22980 10920 23040 10980
rect 23250 10920 23310 10980
rect 23970 10920 24030 10980
rect 24210 10920 24270 10980
rect 25650 10920 25710 10980
rect 25920 10920 25980 10980
rect 26070 10920 26130 10980
rect 26430 10920 26490 10980
rect 26580 10920 26640 10980
rect 26850 10920 26910 10980
rect 28050 10920 28110 10980
rect 28290 10920 28350 10980
rect 29490 10920 29550 10980
rect 30690 10920 30750 10980
rect 31890 10920 31950 10980
rect 32040 10920 32100 10980
rect 32280 10920 32340 10980
rect 33330 10920 33390 10980
rect 33600 10920 33660 10980
rect 33750 10920 33810 10980
rect 34110 10920 34170 10980
rect 34260 10920 34320 10980
rect 34530 10920 34590 10980
rect 35730 10920 35790 10980
rect 35970 10920 36030 10980
rect 36210 10920 36270 10980
rect 36930 10920 36990 10980
rect 37170 10920 37230 10980
rect 37890 10920 37950 10980
rect 38130 10920 38190 10980
rect 38370 10920 38430 10980
rect 39090 10920 39150 10980
rect 39240 10920 39300 10980
rect 39480 10920 39540 10980
rect 40530 10920 40590 10980
rect 40770 10920 40830 10980
rect 41730 10920 41790 10980
rect 41970 10920 42030 10980
rect 42690 10920 42750 10980
rect 42960 10920 43020 10980
rect 43110 10920 43170 10980
rect 43470 10920 43530 10980
rect 43620 10920 43680 10980
rect 43890 10920 43950 10980
rect 45330 10920 45390 10980
rect 45600 10920 45660 10980
rect 45750 10920 45810 10980
rect 46110 10920 46170 10980
rect 46260 10920 46320 10980
rect 46530 10920 46590 10980
rect 47730 10920 47790 10980
rect 47970 10920 48030 10980
rect 49170 10920 49230 10980
rect 49410 10920 49470 10980
rect 5820 10050 5880 10320
rect 5730 8880 5790 9990
rect 6060 9690 6120 9720
rect 5970 9630 6120 9690
rect 5970 9390 6030 9630
rect 6210 9570 6270 9720
rect 6210 9510 6360 9570
rect 5970 9270 6060 9390
rect 5970 8880 6030 9270
rect 6300 9090 6360 9510
rect 6930 9090 6990 10320
rect 6210 8880 6270 9030
rect 6900 8970 6990 9090
rect 7170 9930 7230 10320
rect 7170 9810 7260 9930
rect 7170 8970 7230 9810
rect 7890 9210 7950 9720
rect 8160 9690 8220 9720
rect 8130 9630 8220 9690
rect 8130 9510 8190 9630
rect 6930 8880 6990 8970
rect 7080 8910 7230 8970
rect 7080 8880 7140 8910
rect 7890 8880 7950 9090
rect 8100 8970 8160 9390
rect 8310 9270 8370 9720
rect 8670 9540 8730 9720
rect 8820 9690 8880 9720
rect 9090 9690 9150 9720
rect 8820 9630 9150 9690
rect 8670 9480 8880 9540
rect 8820 9210 8880 9480
rect 9090 9210 9150 9630
rect 8400 9150 8640 9210
rect 8100 8910 8220 8970
rect 8160 8880 8220 8910
rect 8310 8910 8340 9030
rect 8580 8970 8640 9150
rect 9810 9090 9870 10320
rect 10050 9690 10110 10320
rect 10050 9270 10110 9570
rect 10290 9330 10350 10320
rect 11490 9930 11550 10320
rect 11460 9810 11550 9930
rect 10050 9210 10200 9270
rect 9090 8970 9150 9090
rect 9810 9000 9840 9090
rect 8580 8910 8730 8970
rect 8310 8880 8370 8910
rect 8670 8880 8730 8910
rect 8820 8910 9150 8970
rect 8820 8880 8880 8910
rect 9090 8880 9150 8910
rect 9900 8580 9960 8970
rect 10140 8880 10200 9210
rect 10290 9210 10380 9330
rect 10290 8880 10350 9210
rect 11490 8970 11550 9810
rect 11730 9090 11790 10320
rect 13890 9210 13950 9720
rect 14160 9690 14220 9720
rect 14130 9630 14220 9690
rect 14130 9510 14190 9630
rect 11730 8970 11820 9090
rect 11490 8910 11640 8970
rect 11580 8880 11640 8910
rect 11730 8880 11790 8970
rect 13890 8880 13950 9090
rect 14100 8970 14160 9390
rect 14310 9270 14370 9720
rect 14670 9540 14730 9720
rect 14820 9690 14880 9720
rect 15090 9690 15150 9720
rect 14820 9630 15150 9690
rect 14670 9480 14880 9540
rect 14820 9210 14880 9480
rect 15090 9210 15150 9630
rect 14400 9150 14640 9210
rect 14100 8910 14220 8970
rect 14160 8880 14220 8910
rect 14310 8910 14340 9030
rect 14580 8970 14640 9150
rect 16530 9090 16590 10320
rect 15090 8970 15150 9090
rect 16500 8970 16590 9090
rect 16770 9930 16830 10320
rect 16770 9810 16860 9930
rect 16770 8970 16830 9810
rect 21330 9930 21390 10320
rect 21300 9810 21390 9930
rect 17490 9660 17550 9720
rect 17760 9690 17820 9720
rect 17460 9600 17550 9660
rect 17700 9630 17820 9690
rect 17460 9210 17520 9600
rect 17700 9450 17760 9630
rect 17910 9510 17970 9720
rect 14580 8910 14730 8970
rect 14310 8880 14370 8910
rect 14670 8880 14730 8910
rect 14820 8910 15150 8970
rect 14820 8880 14880 8910
rect 15090 8880 15150 8910
rect 16530 8880 16590 8970
rect 16680 8910 16830 8970
rect 16680 8880 16740 8910
rect 17490 8880 17550 9090
rect 17700 8970 17760 9330
rect 18030 9210 18090 9510
rect 18270 9360 18330 9720
rect 18420 9690 18480 9720
rect 18690 9690 18750 9720
rect 18420 9630 18750 9690
rect 18270 9300 18420 9360
rect 18360 9210 18420 9300
rect 18690 9210 18750 9630
rect 19410 9690 19470 9720
rect 19680 9690 19740 9720
rect 19410 9630 19740 9690
rect 19410 9210 19470 9630
rect 19830 9540 19890 9720
rect 19680 9480 19890 9540
rect 19680 9210 19740 9480
rect 20190 9270 20250 9720
rect 20340 9690 20400 9720
rect 20340 9630 20430 9690
rect 20370 9510 20430 9630
rect 18030 9150 18240 9210
rect 17700 8910 17820 8970
rect 17760 8880 17820 8910
rect 17910 8910 17940 8970
rect 18180 8970 18240 9150
rect 19920 9150 20160 9210
rect 18690 8970 18750 9090
rect 18180 8910 18330 8970
rect 17910 8880 17970 8910
rect 18270 8880 18330 8910
rect 18420 8910 18750 8970
rect 18420 8880 18480 8910
rect 18690 8880 18750 8910
rect 19410 8970 19470 9090
rect 19920 8970 19980 9150
rect 19410 8910 19740 8970
rect 19410 8880 19470 8910
rect 19680 8880 19740 8910
rect 19830 8910 19980 8970
rect 20220 8910 20250 9030
rect 20400 8970 20460 9390
rect 20610 9210 20670 9720
rect 19830 8880 19890 8910
rect 20190 8880 20250 8910
rect 20340 8910 20460 8970
rect 20340 8880 20400 8910
rect 20610 8880 20670 9090
rect 21330 8970 21390 9810
rect 21570 9090 21630 10320
rect 22050 9690 22110 9720
rect 22320 9690 22380 9720
rect 22050 9630 22380 9690
rect 22050 9210 22110 9630
rect 22470 9540 22530 9720
rect 22320 9480 22530 9540
rect 22320 9210 22380 9480
rect 22830 9270 22890 9720
rect 22980 9690 23040 9720
rect 22980 9630 23070 9690
rect 23010 9510 23070 9630
rect 22560 9150 22800 9210
rect 21570 8970 21660 9090
rect 22050 8970 22110 9090
rect 22560 8970 22620 9150
rect 21330 8910 21480 8970
rect 21420 8880 21480 8910
rect 21570 8880 21630 8970
rect 22050 8910 22380 8970
rect 22050 8880 22110 8910
rect 22320 8880 22380 8910
rect 22470 8910 22620 8970
rect 22860 8910 22890 9030
rect 23040 8970 23100 9390
rect 23250 9210 23310 9720
rect 23970 9090 24030 10320
rect 22470 8880 22530 8910
rect 22830 8880 22890 8910
rect 22980 8910 23100 8970
rect 22980 8880 23040 8910
rect 23250 8880 23310 9090
rect 23940 8970 24030 9090
rect 24210 9930 24270 10320
rect 24210 9810 24300 9930
rect 24210 8970 24270 9810
rect 25650 9210 25710 9720
rect 25920 9690 25980 9720
rect 25890 9630 25980 9690
rect 25890 9510 25950 9630
rect 23970 8880 24030 8970
rect 24120 8910 24270 8970
rect 24120 8880 24180 8910
rect 25650 8880 25710 9090
rect 25860 8970 25920 9390
rect 26070 9270 26130 9720
rect 26430 9540 26490 9720
rect 26580 9690 26640 9720
rect 26850 9690 26910 9720
rect 26580 9630 26910 9690
rect 26430 9480 26640 9540
rect 26580 9210 26640 9480
rect 26850 9210 26910 9630
rect 26160 9150 26400 9210
rect 25860 8910 25980 8970
rect 25920 8880 25980 8910
rect 26070 8910 26100 9030
rect 26340 8970 26400 9150
rect 28050 9090 28110 10320
rect 26850 8970 26910 9090
rect 28020 8970 28110 9090
rect 28290 9930 28350 10320
rect 28290 9810 28380 9930
rect 28290 8970 28350 9810
rect 26340 8910 26490 8970
rect 26070 8880 26130 8910
rect 26430 8880 26490 8910
rect 26580 8910 26910 8970
rect 26580 8880 26640 8910
rect 26850 8880 26910 8910
rect 28050 8880 28110 8970
rect 28200 8910 28350 8970
rect 28200 8880 28260 8910
rect 29490 8790 29550 10320
rect 30690 8790 30750 10320
rect 32280 10050 32340 10320
rect 31890 9570 31950 9720
rect 32040 9690 32100 9720
rect 32040 9630 32190 9690
rect 31800 9510 31950 9570
rect 31800 9090 31860 9510
rect 32130 9390 32190 9630
rect 32100 9270 32190 9390
rect 31890 8880 31950 9030
rect 32130 8880 32190 9270
rect 32370 8880 32430 9990
rect 33330 9690 33390 9720
rect 33600 9690 33660 9720
rect 33330 9630 33660 9690
rect 33330 9210 33390 9630
rect 33750 9360 33810 9720
rect 33660 9300 33810 9360
rect 34110 9510 34170 9720
rect 34260 9690 34320 9720
rect 34260 9630 34380 9690
rect 33660 9210 33720 9300
rect 33990 9210 34050 9510
rect 33840 9150 34050 9210
rect 34320 9450 34380 9630
rect 34530 9660 34590 9720
rect 34530 9600 34620 9660
rect 33330 8970 33390 9090
rect 33840 8970 33900 9150
rect 33330 8910 33660 8970
rect 33330 8880 33390 8910
rect 33600 8880 33660 8910
rect 33750 8910 33900 8970
rect 34320 8970 34380 9330
rect 34560 9210 34620 9600
rect 35730 9090 35790 10320
rect 35970 9690 36030 10320
rect 35970 9270 36030 9570
rect 36210 9330 36270 10320
rect 35970 9210 36120 9270
rect 34140 8910 34170 8970
rect 33750 8880 33810 8910
rect 34110 8880 34170 8910
rect 34260 8910 34380 8970
rect 34260 8880 34320 8910
rect 34530 8880 34590 9090
rect 35730 9000 35760 9090
rect 29490 8670 29580 8790
rect 30660 8670 30750 8790
rect 29490 8580 29550 8670
rect 30690 8580 30750 8670
rect 35820 8580 35880 8970
rect 36060 8880 36120 9210
rect 36210 9210 36300 9330
rect 36210 8880 36270 9210
rect 36930 9090 36990 10320
rect 36900 8970 36990 9090
rect 37170 9930 37230 10320
rect 37170 9810 37260 9930
rect 37170 8970 37230 9810
rect 37890 9090 37950 10320
rect 38130 9690 38190 10320
rect 38130 9270 38190 9570
rect 38370 9330 38430 10320
rect 39480 10050 39540 10320
rect 39090 9570 39150 9720
rect 39240 9690 39300 9720
rect 39240 9630 39390 9690
rect 39000 9510 39150 9570
rect 38130 9210 38280 9270
rect 37890 9000 37920 9090
rect 36930 8880 36990 8970
rect 37080 8910 37230 8970
rect 37080 8880 37140 8910
rect 37980 8580 38040 8970
rect 38220 8880 38280 9210
rect 38370 9210 38460 9330
rect 38370 8880 38430 9210
rect 39000 9090 39060 9510
rect 39330 9390 39390 9630
rect 39300 9270 39390 9390
rect 39090 8880 39150 9030
rect 39330 8880 39390 9270
rect 39570 8880 39630 9990
rect 40530 9090 40590 10320
rect 40500 8970 40590 9090
rect 40770 9930 40830 10320
rect 40770 9810 40860 9930
rect 40770 8970 40830 9810
rect 41730 9090 41790 10320
rect 41700 8970 41790 9090
rect 41970 9930 42030 10320
rect 41970 9810 42060 9930
rect 41970 8970 42030 9810
rect 47730 9930 47790 10320
rect 47700 9810 47790 9930
rect 42690 9210 42750 9720
rect 42960 9690 43020 9720
rect 42930 9630 43020 9690
rect 42930 9510 42990 9630
rect 40530 8880 40590 8970
rect 40680 8910 40830 8970
rect 40680 8880 40740 8910
rect 41730 8880 41790 8970
rect 41880 8910 42030 8970
rect 41880 8880 41940 8910
rect 42690 8880 42750 9090
rect 42900 8970 42960 9390
rect 43110 9270 43170 9720
rect 43470 9540 43530 9720
rect 43620 9690 43680 9720
rect 43890 9690 43950 9720
rect 43620 9630 43950 9690
rect 43470 9480 43680 9540
rect 43620 9210 43680 9480
rect 43890 9210 43950 9630
rect 45330 9210 45390 9720
rect 45600 9690 45660 9720
rect 45570 9630 45660 9690
rect 45570 9510 45630 9630
rect 43200 9150 43440 9210
rect 42900 8910 43020 8970
rect 42960 8880 43020 8910
rect 43110 8910 43140 9030
rect 43380 8970 43440 9150
rect 43890 8970 43950 9090
rect 43380 8910 43530 8970
rect 43110 8880 43170 8910
rect 43470 8880 43530 8910
rect 43620 8910 43950 8970
rect 43620 8880 43680 8910
rect 43890 8880 43950 8910
rect 45330 8880 45390 9090
rect 45540 8970 45600 9390
rect 45750 9270 45810 9720
rect 46110 9540 46170 9720
rect 46260 9690 46320 9720
rect 46530 9690 46590 9720
rect 46260 9630 46590 9690
rect 46110 9480 46320 9540
rect 46260 9210 46320 9480
rect 46530 9210 46590 9630
rect 45840 9150 46080 9210
rect 45540 8910 45660 8970
rect 45600 8880 45660 8910
rect 45750 8910 45780 9030
rect 46020 8970 46080 9150
rect 46530 8970 46590 9090
rect 46020 8910 46170 8970
rect 45750 8880 45810 8910
rect 46110 8880 46170 8910
rect 46260 8910 46590 8970
rect 47730 8970 47790 9810
rect 47970 9090 48030 10320
rect 49170 9930 49230 10320
rect 49140 9810 49230 9930
rect 47970 8970 48060 9090
rect 49170 8970 49230 9810
rect 49410 9090 49470 10320
rect 49410 8970 49500 9090
rect 47730 8910 47880 8970
rect 46260 8880 46320 8910
rect 46530 8880 46590 8910
rect 47820 8880 47880 8910
rect 47970 8880 48030 8970
rect 49170 8910 49320 8970
rect 49260 8880 49320 8910
rect 49410 8880 49470 8970
rect 5730 8220 5790 8280
rect 5970 8220 6030 8280
rect 6210 8220 6270 8280
rect 6930 8220 6990 8280
rect 7080 8220 7140 8280
rect 7890 8220 7950 8280
rect 8160 8220 8220 8280
rect 8310 8220 8370 8280
rect 8670 8220 8730 8280
rect 8820 8220 8880 8280
rect 9090 8220 9150 8280
rect 9900 8220 9960 8280
rect 10140 8220 10200 8280
rect 10290 8220 10350 8280
rect 11580 8220 11640 8280
rect 11730 8220 11790 8280
rect 13890 8220 13950 8280
rect 14160 8220 14220 8280
rect 14310 8220 14370 8280
rect 14670 8220 14730 8280
rect 14820 8220 14880 8280
rect 15090 8220 15150 8280
rect 16530 8220 16590 8280
rect 16680 8220 16740 8280
rect 17490 8220 17550 8280
rect 17760 8220 17820 8280
rect 17910 8220 17970 8280
rect 18270 8220 18330 8280
rect 18420 8220 18480 8280
rect 18690 8220 18750 8280
rect 19410 8220 19470 8280
rect 19680 8220 19740 8280
rect 19830 8220 19890 8280
rect 20190 8220 20250 8280
rect 20340 8220 20400 8280
rect 20610 8220 20670 8280
rect 21420 8220 21480 8280
rect 21570 8220 21630 8280
rect 22050 8220 22110 8280
rect 22320 8220 22380 8280
rect 22470 8220 22530 8280
rect 22830 8220 22890 8280
rect 22980 8220 23040 8280
rect 23250 8220 23310 8280
rect 23970 8220 24030 8280
rect 24120 8220 24180 8280
rect 25650 8220 25710 8280
rect 25920 8220 25980 8280
rect 26070 8220 26130 8280
rect 26430 8220 26490 8280
rect 26580 8220 26640 8280
rect 26850 8220 26910 8280
rect 28050 8220 28110 8280
rect 28200 8220 28260 8280
rect 29490 8220 29550 8280
rect 30690 8220 30750 8280
rect 31890 8220 31950 8280
rect 32130 8220 32190 8280
rect 32370 8220 32430 8280
rect 33330 8220 33390 8280
rect 33600 8220 33660 8280
rect 33750 8220 33810 8280
rect 34110 8220 34170 8280
rect 34260 8220 34320 8280
rect 34530 8220 34590 8280
rect 35820 8220 35880 8280
rect 36060 8220 36120 8280
rect 36210 8220 36270 8280
rect 36930 8220 36990 8280
rect 37080 8220 37140 8280
rect 37980 8220 38040 8280
rect 38220 8220 38280 8280
rect 38370 8220 38430 8280
rect 39090 8220 39150 8280
rect 39330 8220 39390 8280
rect 39570 8220 39630 8280
rect 40530 8220 40590 8280
rect 40680 8220 40740 8280
rect 41730 8220 41790 8280
rect 41880 8220 41940 8280
rect 42690 8220 42750 8280
rect 42960 8220 43020 8280
rect 43110 8220 43170 8280
rect 43470 8220 43530 8280
rect 43620 8220 43680 8280
rect 43890 8220 43950 8280
rect 45330 8220 45390 8280
rect 45600 8220 45660 8280
rect 45750 8220 45810 8280
rect 46110 8220 46170 8280
rect 46260 8220 46320 8280
rect 46530 8220 46590 8280
rect 47820 8220 47880 8280
rect 47970 8220 48030 8280
rect 49260 8220 49320 8280
rect 49410 8220 49470 8280
rect 5730 7920 5790 7980
rect 6000 7920 6060 7980
rect 6150 7920 6210 7980
rect 6510 7920 6570 7980
rect 6660 7920 6720 7980
rect 6930 7920 6990 7980
rect 8130 7920 8190 7980
rect 8850 7920 8910 7980
rect 9090 7920 9150 7980
rect 9330 7920 9390 7980
rect 10050 7920 10110 7980
rect 10200 7920 10260 7980
rect 11010 7920 11070 7980
rect 11250 7920 11310 7980
rect 11490 7920 11550 7980
rect 12450 7920 12510 7980
rect 12600 7920 12660 7980
rect 13980 7920 14040 7980
rect 14130 7920 14190 7980
rect 14370 7920 14430 7980
rect 15570 7920 15630 7980
rect 15810 7920 15870 7980
rect 18210 7920 18270 7980
rect 18450 7920 18510 7980
rect 20850 7920 20910 7980
rect 21000 7920 21060 7980
rect 23490 7920 23550 7980
rect 23640 7920 23700 7980
rect 25890 7920 25950 7980
rect 26160 7920 26220 7980
rect 26310 7920 26370 7980
rect 26670 7920 26730 7980
rect 26820 7920 26880 7980
rect 27090 7920 27150 7980
rect 28050 7920 28110 7980
rect 28200 7920 28260 7980
rect 29250 7920 29310 7980
rect 29400 7920 29460 7980
rect 30210 7920 30270 7980
rect 30480 7920 30540 7980
rect 30630 7920 30690 7980
rect 30990 7920 31050 7980
rect 31140 7920 31200 7980
rect 31410 7920 31470 7980
rect 32130 7920 32190 7980
rect 32370 7920 32430 7980
rect 32610 7920 32670 7980
rect 33330 7920 33390 7980
rect 33480 7920 33540 7980
rect 34860 7920 34920 7980
rect 35010 7920 35070 7980
rect 36210 7920 36270 7980
rect 36360 7920 36420 7980
rect 37650 7920 37710 7980
rect 37890 7920 37950 7980
rect 38130 7920 38190 7980
rect 39090 7920 39150 7980
rect 39240 7920 39300 7980
rect 40530 7920 40590 7980
rect 40680 7920 40740 7980
rect 43410 7920 43470 7980
rect 43650 7920 43710 7980
rect 44670 7920 44730 7980
rect 44820 7920 44880 7980
rect 45180 7920 45240 7980
rect 45330 7920 45390 7980
rect 46530 7920 46590 7980
rect 47490 7920 47550 7980
rect 47730 7920 47790 7980
rect 47970 7920 48030 7980
rect 8130 7530 8190 7620
rect 8130 7410 8220 7530
rect 5730 7290 5790 7320
rect 6000 7290 6060 7320
rect 5730 7230 6060 7290
rect 6150 7290 6210 7320
rect 6510 7290 6570 7320
rect 6150 7230 6300 7290
rect 5730 7110 5790 7230
rect 6240 7050 6300 7230
rect 6540 7170 6570 7290
rect 6660 7290 6720 7320
rect 6660 7230 6780 7290
rect 6240 6990 6480 7050
rect 5730 6570 5790 6990
rect 6000 6720 6060 6990
rect 6000 6660 6210 6720
rect 5730 6510 6060 6570
rect 5730 6480 5790 6510
rect 6000 6480 6060 6510
rect 6150 6480 6210 6660
rect 6510 6480 6570 6930
rect 6720 6810 6780 7230
rect 6930 7110 6990 7320
rect 6690 6570 6750 6690
rect 6660 6510 6750 6570
rect 6660 6480 6720 6510
rect 6930 6480 6990 6990
rect 8130 5880 8190 7410
rect 8850 6210 8910 7320
rect 9090 6930 9150 7320
rect 9330 7170 9390 7320
rect 10050 7230 10110 7320
rect 10200 7290 10260 7320
rect 10200 7230 10350 7290
rect 10020 7110 10110 7230
rect 9090 6810 9180 6930
rect 9090 6570 9150 6810
rect 9420 6690 9480 7110
rect 9330 6630 9480 6690
rect 9090 6510 9240 6570
rect 9180 6480 9240 6510
rect 9330 6480 9390 6630
rect 8940 5880 9000 6150
rect 10050 5880 10110 7110
rect 10290 6390 10350 7230
rect 10290 6270 10380 6390
rect 10290 5880 10350 6270
rect 11010 6210 11070 7320
rect 11250 6930 11310 7320
rect 11490 7170 11550 7320
rect 12450 7230 12510 7320
rect 12600 7290 12660 7320
rect 13980 7290 14040 7320
rect 12600 7230 12750 7290
rect 12420 7110 12510 7230
rect 11250 6810 11340 6930
rect 11250 6570 11310 6810
rect 11580 6690 11640 7110
rect 11490 6630 11640 6690
rect 11250 6510 11400 6570
rect 11340 6480 11400 6510
rect 11490 6480 11550 6630
rect 11100 5880 11160 6150
rect 12450 5880 12510 7110
rect 12690 6390 12750 7230
rect 13800 7230 14040 7290
rect 13800 6690 13860 7230
rect 14130 6990 14190 7320
rect 14100 6870 14190 6990
rect 13890 6480 13950 6630
rect 14130 6480 14190 6870
rect 14370 6480 14430 7620
rect 15570 7530 15630 7620
rect 15540 7410 15630 7530
rect 15570 6480 15630 7410
rect 15810 6690 15870 7620
rect 18210 7530 18270 7620
rect 18180 7410 18270 7530
rect 15810 6570 15900 6690
rect 15720 6510 15870 6570
rect 15720 6480 15780 6510
rect 18210 6480 18270 7410
rect 18450 6690 18510 7620
rect 43410 7530 43470 7620
rect 43380 7410 43470 7530
rect 20850 7230 20910 7320
rect 21000 7290 21060 7320
rect 21000 7230 21150 7290
rect 23490 7230 23550 7320
rect 23640 7290 23700 7320
rect 23640 7230 23790 7290
rect 20820 7110 20910 7230
rect 18450 6570 18540 6690
rect 18360 6510 18510 6570
rect 18360 6480 18420 6510
rect 12690 6270 12780 6390
rect 12690 5880 12750 6270
rect 20850 5880 20910 7110
rect 21090 6390 21150 7230
rect 23460 7110 23550 7230
rect 21090 6270 21180 6390
rect 21090 5880 21150 6270
rect 23490 5880 23550 7110
rect 23730 6390 23790 7230
rect 25890 7110 25950 7320
rect 26160 7290 26220 7320
rect 26100 7230 26220 7290
rect 26310 7290 26370 7320
rect 26670 7290 26730 7320
rect 26310 7230 26340 7290
rect 25860 6600 25920 6990
rect 26100 6870 26160 7230
rect 26580 7230 26730 7290
rect 26820 7290 26880 7320
rect 27090 7290 27150 7320
rect 26820 7230 27150 7290
rect 28050 7230 28110 7320
rect 28200 7290 28260 7320
rect 28200 7230 28350 7290
rect 29250 7230 29310 7320
rect 29400 7290 29460 7320
rect 29400 7230 29550 7290
rect 26580 7050 26640 7230
rect 27090 7110 27150 7230
rect 28020 7110 28110 7230
rect 25860 6540 25950 6600
rect 25890 6480 25950 6540
rect 26100 6570 26160 6750
rect 26430 6990 26640 7050
rect 26430 6690 26490 6990
rect 26760 6900 26820 6990
rect 26100 6510 26220 6570
rect 26160 6480 26220 6510
rect 26310 6480 26370 6690
rect 26670 6840 26820 6900
rect 26670 6480 26730 6840
rect 27090 6570 27150 6990
rect 26820 6510 27150 6570
rect 26820 6480 26880 6510
rect 27090 6480 27150 6510
rect 23730 6270 23820 6390
rect 23730 5880 23790 6270
rect 28050 5880 28110 7110
rect 28290 6390 28350 7230
rect 29220 7110 29310 7230
rect 28290 6270 28380 6390
rect 28290 5880 28350 6270
rect 29250 5880 29310 7110
rect 29490 6390 29550 7230
rect 30210 7110 30270 7320
rect 30480 7290 30540 7320
rect 30420 7230 30540 7290
rect 30630 7290 30690 7320
rect 30990 7290 31050 7320
rect 30210 6480 30270 6990
rect 30420 6810 30480 7230
rect 30630 7170 30660 7290
rect 30900 7230 31050 7290
rect 31140 7290 31200 7320
rect 31410 7290 31470 7320
rect 31140 7230 31470 7290
rect 30900 7050 30960 7230
rect 31410 7110 31470 7230
rect 32130 7170 32190 7320
rect 30720 6990 30960 7050
rect 30450 6570 30510 6690
rect 30450 6510 30540 6570
rect 30480 6480 30540 6510
rect 30630 6480 30690 6930
rect 31140 6720 31200 6990
rect 30990 6660 31200 6720
rect 30990 6480 31050 6660
rect 31410 6570 31470 6990
rect 32040 6690 32100 7110
rect 32370 6930 32430 7320
rect 32340 6810 32430 6930
rect 32040 6630 32190 6690
rect 31140 6510 31470 6570
rect 31140 6480 31200 6510
rect 31410 6480 31470 6510
rect 32130 6480 32190 6630
rect 32370 6570 32430 6810
rect 32280 6510 32430 6570
rect 32280 6480 32340 6510
rect 29490 6270 29580 6390
rect 29490 5880 29550 6270
rect 32610 6210 32670 7320
rect 33330 7230 33390 7320
rect 33480 7290 33540 7320
rect 34860 7290 34920 7320
rect 33480 7230 33630 7290
rect 33300 7110 33390 7230
rect 32520 5880 32580 6150
rect 33330 5880 33390 7110
rect 33570 6390 33630 7230
rect 34770 7230 34920 7290
rect 35010 7230 35070 7320
rect 36210 7230 36270 7320
rect 36360 7290 36420 7320
rect 36360 7230 36510 7290
rect 34770 6390 34830 7230
rect 33570 6270 33660 6390
rect 34740 6270 34830 6390
rect 33570 5880 33630 6270
rect 34770 5880 34830 6270
rect 35010 7110 35100 7230
rect 36180 7110 36270 7230
rect 35010 5880 35070 7110
rect 36210 5880 36270 7110
rect 36450 6390 36510 7230
rect 36450 6270 36540 6390
rect 36450 5880 36510 6270
rect 37650 6210 37710 7320
rect 37890 6930 37950 7320
rect 38130 7170 38190 7320
rect 39090 7230 39150 7320
rect 39240 7290 39300 7320
rect 39240 7230 39390 7290
rect 40530 7230 40590 7320
rect 40680 7290 40740 7320
rect 40680 7230 40830 7290
rect 39060 7110 39150 7230
rect 37890 6810 37980 6930
rect 37890 6570 37950 6810
rect 38220 6690 38280 7110
rect 38130 6630 38280 6690
rect 37890 6510 38040 6570
rect 37980 6480 38040 6510
rect 38130 6480 38190 6630
rect 37740 5880 37800 6150
rect 39090 5880 39150 7110
rect 39330 6390 39390 7230
rect 40500 7110 40590 7230
rect 39330 6270 39420 6390
rect 39330 5880 39390 6270
rect 40530 5880 40590 7110
rect 40770 6390 40830 7230
rect 43410 6480 43470 7410
rect 43650 6690 43710 7620
rect 46530 7530 46590 7620
rect 46530 7410 46620 7530
rect 44670 7290 44730 7320
rect 44520 7230 44730 7290
rect 44520 6690 44580 7230
rect 43650 6570 43740 6690
rect 43560 6510 43710 6570
rect 43560 6480 43620 6510
rect 44610 6480 44670 6630
rect 44820 6570 44880 7320
rect 45180 7290 45240 7320
rect 45120 7230 45240 7290
rect 45330 7230 45390 7320
rect 45120 6930 45180 7230
rect 45330 7170 45450 7230
rect 45120 6900 45150 6930
rect 44820 6510 44910 6570
rect 44850 6480 44910 6510
rect 45090 6480 45150 6900
rect 45390 6690 45450 7170
rect 45390 6570 45420 6690
rect 45330 6510 45450 6570
rect 45330 6480 45390 6510
rect 40770 6270 40860 6390
rect 40770 5880 40830 6270
rect 46530 5880 46590 7410
rect 47490 6210 47550 7320
rect 47730 6930 47790 7320
rect 47970 7170 48030 7320
rect 47730 6810 47820 6930
rect 47730 6570 47790 6810
rect 48060 6690 48120 7110
rect 47970 6630 48120 6690
rect 47730 6510 47880 6570
rect 47820 6480 47880 6510
rect 47970 6480 48030 6630
rect 47580 5880 47640 6150
rect 5730 5220 5790 5280
rect 6000 5220 6060 5280
rect 6150 5220 6210 5280
rect 6510 5220 6570 5280
rect 6660 5220 6720 5280
rect 6930 5220 6990 5280
rect 8130 5220 8190 5280
rect 8940 5220 9000 5280
rect 9180 5220 9240 5280
rect 9330 5220 9390 5280
rect 10050 5220 10110 5280
rect 10290 5220 10350 5280
rect 11100 5220 11160 5280
rect 11340 5220 11400 5280
rect 11490 5220 11550 5280
rect 12450 5220 12510 5280
rect 12690 5220 12750 5280
rect 13890 5220 13950 5280
rect 14130 5220 14190 5280
rect 14370 5220 14430 5280
rect 15570 5220 15630 5280
rect 15720 5220 15780 5280
rect 18210 5220 18270 5280
rect 18360 5220 18420 5280
rect 20850 5220 20910 5280
rect 21090 5220 21150 5280
rect 23490 5220 23550 5280
rect 23730 5220 23790 5280
rect 25890 5220 25950 5280
rect 26160 5220 26220 5280
rect 26310 5220 26370 5280
rect 26670 5220 26730 5280
rect 26820 5220 26880 5280
rect 27090 5220 27150 5280
rect 28050 5220 28110 5280
rect 28290 5220 28350 5280
rect 29250 5220 29310 5280
rect 29490 5220 29550 5280
rect 30210 5220 30270 5280
rect 30480 5220 30540 5280
rect 30630 5220 30690 5280
rect 30990 5220 31050 5280
rect 31140 5220 31200 5280
rect 31410 5220 31470 5280
rect 32130 5220 32190 5280
rect 32280 5220 32340 5280
rect 32520 5220 32580 5280
rect 33330 5220 33390 5280
rect 33570 5220 33630 5280
rect 34770 5220 34830 5280
rect 35010 5220 35070 5280
rect 36210 5220 36270 5280
rect 36450 5220 36510 5280
rect 37740 5220 37800 5280
rect 37980 5220 38040 5280
rect 38130 5220 38190 5280
rect 39090 5220 39150 5280
rect 39330 5220 39390 5280
rect 40530 5220 40590 5280
rect 40770 5220 40830 5280
rect 43410 5220 43470 5280
rect 43560 5220 43620 5280
rect 44610 5220 44670 5280
rect 44850 5220 44910 5280
rect 45090 5220 45150 5280
rect 45330 5220 45390 5280
rect 46530 5220 46590 5280
rect 47580 5220 47640 5280
rect 47820 5220 47880 5280
rect 47970 5220 48030 5280
<< polycontact >>
rect 6180 43050 6300 43170
rect 6780 43110 6900 43230
rect 6060 42810 6180 42930
rect 5700 42090 5820 42210
rect 7260 42270 7380 42390
rect 8340 43050 8460 43170
rect 8220 42810 8340 42930
rect 9060 42990 9180 43110
rect 9540 43170 9660 43290
rect 9480 42930 9600 43050
rect 9960 42990 10080 43110
rect 10260 42990 10380 43110
rect 9270 42690 9390 42810
rect 10860 42570 10980 42690
rect 11340 43410 11460 43530
rect 12300 42570 12420 42690
rect 12780 43410 12900 43530
rect 21180 43410 21300 43530
rect 13860 43050 13980 43170
rect 13980 42810 14100 42930
rect 7860 42090 7980 42210
rect 15420 43110 15540 43230
rect 14340 42090 14460 42210
rect 17220 43050 17340 43170
rect 17340 42810 17460 42930
rect 15900 42270 16020 42390
rect 19380 42990 19500 43110
rect 19680 42990 19800 43110
rect 20100 43170 20220 43290
rect 20580 42990 20700 43110
rect 20400 42750 20520 42870
rect 20070 42570 20190 42690
rect 17700 42090 17820 42210
rect 34620 43410 34740 43530
rect 22740 42990 22860 43110
rect 23220 43170 23340 43290
rect 23160 42930 23280 43050
rect 23640 42990 23760 43110
rect 23940 42990 24060 43110
rect 22950 42690 23070 42810
rect 25620 43050 25740 43170
rect 26700 43110 26820 43230
rect 25500 42810 25620 42930
rect 25140 42090 25260 42210
rect 28020 43050 28140 43170
rect 28140 42810 28260 42930
rect 27180 42270 27300 42390
rect 29100 43110 29220 43230
rect 28500 42090 28620 42210
rect 30420 43050 30540 43170
rect 30540 42810 30660 42930
rect 29580 42270 29700 42390
rect 31860 43050 31980 43170
rect 31980 42810 32100 42930
rect 30900 42090 31020 42210
rect 33180 42270 33300 42390
rect 32340 42090 32460 42210
rect 33660 43110 33780 43230
rect 41820 43410 41940 43530
rect 35940 42990 36060 43110
rect 35100 42570 35220 42690
rect 36420 43170 36540 43290
rect 36360 42930 36480 43050
rect 36840 42990 36960 43110
rect 37140 42990 37260 43110
rect 36150 42690 36270 42810
rect 38340 43050 38460 43170
rect 38220 42810 38340 42930
rect 39540 42990 39660 43110
rect 39840 42990 39960 43110
rect 40260 43170 40380 43290
rect 40320 42930 40440 43050
rect 40740 42990 40860 43110
rect 40530 42690 40650 42810
rect 37860 42090 37980 42210
rect 45420 43410 45540 43530
rect 43140 43050 43260 43170
rect 43260 42810 43380 42930
rect 44340 43050 44460 43170
rect 44460 42810 44580 42930
rect 43620 42090 43740 42210
rect 44820 42090 44940 42210
rect 45780 42990 45900 43110
rect 46260 43170 46380 43290
rect 46200 42930 46320 43050
rect 46680 42990 46800 43110
rect 46980 42990 47100 43110
rect 47460 42990 47580 43110
rect 45990 42690 46110 42810
rect 47940 43170 48060 43290
rect 47880 42930 48000 43050
rect 48360 42990 48480 43110
rect 48660 42990 48780 43110
rect 47670 42690 47790 42810
rect 8220 39810 8340 39930
rect 5940 39450 6060 39570
rect 6060 39210 6180 39330
rect 8700 38970 8820 39090
rect 9660 38970 9780 39090
rect 10140 39810 10260 39930
rect 6510 38670 6630 38790
rect 10650 38670 10770 38790
rect 11220 39450 11340 39570
rect 11100 39210 11220 39330
rect 12210 39510 12330 39630
rect 11880 39330 12000 39450
rect 11700 39090 11820 39210
rect 12180 38910 12300 39030
rect 12600 39090 12720 39210
rect 12900 39090 13020 39210
rect 13500 38970 13620 39090
rect 13980 39810 14100 39930
rect 14850 39570 14970 39690
rect 14640 38970 14760 39090
rect 15180 39210 15300 39330
rect 16980 39990 17100 40110
rect 17700 39990 17820 40110
rect 16620 39270 16740 39390
rect 16500 39030 16620 39150
rect 18060 39270 18180 39390
rect 18180 39030 18300 39150
rect 15660 38670 15780 38790
rect 19860 39990 19980 40110
rect 19500 39270 19620 39390
rect 19380 39030 19500 39150
rect 20940 39810 21060 39930
rect 25380 39990 25500 40110
rect 22230 39390 22350 39510
rect 22020 39090 22140 39210
rect 21420 38970 21540 39090
rect 22440 39150 22560 39270
rect 22500 38910 22620 39030
rect 22920 39090 23040 39210
rect 23220 39090 23340 39210
rect 18780 38670 18900 38790
rect 23820 38670 23940 38790
rect 24300 39510 24420 39630
rect 25020 39270 25140 39390
rect 24900 39030 25020 39150
rect 26340 39450 26460 39570
rect 26460 39210 26580 39330
rect 27180 39510 27300 39630
rect 26910 39270 27030 39390
rect 30540 39810 30660 39930
rect 31980 39810 32100 39930
rect 31020 38970 31140 39090
rect 36660 39990 36780 40110
rect 33750 39390 33870 39510
rect 33540 39090 33660 39210
rect 32460 38970 32580 39090
rect 33960 39150 34080 39270
rect 34020 38910 34140 39030
rect 34440 39090 34560 39210
rect 34740 39090 34860 39210
rect 36300 39270 36420 39390
rect 36180 39030 36300 39150
rect 37740 39810 37860 39930
rect 39540 39990 39660 40110
rect 39180 39270 39300 39390
rect 38220 38970 38340 39090
rect 39060 39030 39180 39150
rect 40380 38970 40500 39090
rect 40860 39810 40980 39930
rect 28140 38670 28260 38790
rect 43620 39990 43740 40110
rect 43260 39270 43380 39390
rect 43140 39030 43260 39150
rect 41820 38670 41940 38790
rect 46020 39990 46140 40110
rect 48180 39990 48300 40110
rect 46380 39270 46500 39390
rect 46500 39030 46620 39150
rect 47820 39270 47940 39390
rect 47700 39030 47820 39150
rect 49260 39810 49380 39930
rect 49740 38970 49860 39090
rect 44700 38670 44820 38790
rect 7260 37410 7380 37530
rect 5580 36270 5700 36390
rect 6060 37110 6180 37230
rect 8820 37050 8940 37170
rect 10860 37110 10980 37230
rect 8700 36810 8820 36930
rect 8340 36090 8460 36210
rect 11340 36270 11460 36390
rect 12660 37050 12780 37170
rect 12540 36810 12660 36930
rect 12180 36090 12300 36210
rect 23820 37410 23940 37530
rect 15540 37050 15660 37170
rect 16800 37110 16920 37230
rect 15420 36810 15540 36930
rect 15060 36090 15180 36210
rect 18060 37110 18180 37230
rect 17340 36870 17460 36990
rect 17010 36510 17130 36630
rect 19500 37110 19620 37230
rect 18540 36270 18660 36390
rect 20940 37110 21060 37230
rect 19980 36270 20100 36390
rect 22380 37110 22500 37230
rect 21420 36270 21540 36390
rect 22860 36270 22980 36390
rect 31260 37410 31380 37530
rect 25020 36270 25140 36390
rect 25500 37110 25620 37230
rect 26580 37050 26700 37170
rect 26700 36810 26820 36930
rect 27900 37110 28020 37230
rect 27060 36090 27180 36210
rect 29100 37110 29220 37230
rect 28380 36270 28500 36390
rect 30180 37050 30300 37170
rect 30300 36810 30420 36930
rect 29580 36270 29700 36390
rect 30660 36090 30780 36210
rect 38940 37410 39060 37530
rect 32580 37050 32700 37170
rect 32460 36810 32580 36930
rect 32100 36090 32220 36210
rect 33180 36270 33300 36390
rect 33660 37110 33780 37230
rect 34620 37110 34740 37230
rect 35700 36990 35820 37110
rect 36000 36990 36120 37110
rect 36420 37170 36540 37290
rect 36480 36930 36600 37050
rect 36900 36990 37020 37110
rect 36690 36690 36810 36810
rect 35100 36270 35220 36390
rect 41580 37410 41700 37530
rect 40170 36810 40290 36930
rect 39900 36570 40020 36690
rect 40620 36870 40740 36990
rect 40740 36630 40860 36750
rect 43740 37410 43860 37530
rect 42900 37050 43020 37170
rect 42780 36810 42900 36930
rect 42420 36090 42540 36210
rect 44580 37050 44700 37170
rect 44700 36810 44820 36930
rect 46140 37110 46260 37230
rect 45060 36090 45180 36210
rect 47700 37050 47820 37170
rect 47820 36810 47940 36930
rect 46620 36270 46740 36390
rect 49260 36270 49380 36390
rect 48180 36090 48300 36210
rect 49740 37110 49860 37230
rect 6660 33990 6780 34110
rect 7860 33990 7980 34110
rect 7020 33270 7140 33390
rect 7140 33030 7260 33150
rect 8220 33270 8340 33390
rect 8340 33030 8460 33150
rect 9570 33510 9690 33630
rect 9240 33330 9360 33450
rect 9060 33090 9180 33210
rect 11730 33510 11850 33630
rect 11400 33330 11520 33450
rect 9540 32910 9660 33030
rect 9960 33090 10080 33210
rect 10260 33090 10380 33210
rect 11220 33090 11340 33210
rect 11700 32910 11820 33030
rect 12120 33090 12240 33210
rect 12420 33090 12540 33210
rect 15180 32970 15300 33090
rect 15660 33810 15780 33930
rect 17220 33990 17340 34110
rect 16860 33270 16980 33390
rect 16740 33030 16860 33150
rect 19260 33810 19380 33930
rect 21090 33570 21210 33690
rect 23940 33990 24060 34110
rect 19740 32970 19860 33090
rect 20880 32970 21000 33090
rect 13980 32670 14100 32790
rect 21420 33210 21540 33330
rect 23580 33270 23700 33390
rect 23460 33030 23580 33150
rect 25380 33990 25500 34110
rect 25020 33270 25140 33390
rect 24900 33030 25020 33150
rect 26310 33390 26430 33510
rect 26100 33090 26220 33210
rect 26520 33150 26640 33270
rect 26580 32910 26700 33030
rect 27000 33090 27120 33210
rect 27300 33090 27420 33210
rect 31020 33810 31140 33930
rect 32580 33990 32700 34110
rect 32220 33270 32340 33390
rect 31500 32970 31620 33090
rect 32100 33030 32220 33150
rect 33180 32970 33300 33090
rect 33660 33810 33780 33930
rect 34620 32970 34740 33090
rect 35100 33810 35220 33930
rect 36060 32970 36180 33090
rect 36540 33810 36660 33930
rect 37500 33810 37620 33930
rect 37980 32970 38100 33090
rect 38940 32970 39060 33090
rect 39420 33810 39540 33930
rect 40740 33990 40860 34110
rect 40380 33270 40500 33390
rect 40260 33030 40380 33150
rect 41580 32970 41700 33090
rect 42060 33810 42180 33930
rect 43620 33990 43740 34110
rect 43260 33270 43380 33390
rect 43140 33030 43260 33150
rect 46740 33990 46860 34110
rect 44550 33390 44670 33510
rect 44340 33090 44460 33210
rect 44760 33150 44880 33270
rect 44820 32910 44940 33030
rect 45240 33090 45360 33210
rect 45540 33090 45660 33210
rect 46380 33270 46500 33390
rect 46260 33030 46380 33150
rect 47580 33810 47700 33930
rect 49020 33810 49140 33930
rect 48060 32970 48180 33090
rect 49500 32970 49620 33090
rect 30540 32670 30660 32790
rect 24060 31410 24180 31530
rect 5460 30990 5580 31110
rect 5760 30990 5880 31110
rect 6180 31170 6300 31290
rect 6660 30990 6780 31110
rect 6480 30750 6600 30870
rect 6150 30570 6270 30690
rect 8100 31050 8220 31170
rect 8220 30810 8340 30930
rect 9660 30270 9780 30390
rect 8580 30090 8700 30210
rect 10140 31110 10260 31230
rect 11220 30990 11340 31110
rect 11700 31170 11820 31290
rect 11640 30930 11760 31050
rect 12120 30990 12240 31110
rect 12420 30990 12540 31110
rect 14820 30990 14940 31110
rect 11430 30690 11550 30810
rect 15300 31170 15420 31290
rect 15000 30750 15120 30870
rect 15720 30990 15840 31110
rect 16020 30990 16140 31110
rect 17220 30990 17340 31110
rect 15330 30570 15450 30690
rect 17700 31170 17820 31290
rect 17400 30750 17520 30870
rect 18120 30990 18240 31110
rect 18420 30990 18540 31110
rect 19380 30990 19500 31110
rect 17730 30570 17850 30690
rect 19860 31170 19980 31290
rect 21180 31110 21300 31230
rect 19800 30930 19920 31050
rect 20280 30990 20400 31110
rect 20580 30990 20700 31110
rect 19590 30690 19710 30810
rect 21660 30270 21780 30390
rect 22740 31050 22860 31170
rect 22620 30810 22740 30930
rect 22260 30090 22380 30210
rect 27420 31410 27540 31530
rect 24960 31110 25080 31230
rect 25500 30870 25620 30990
rect 25170 30510 25290 30630
rect 26580 31050 26700 31170
rect 26460 30810 26580 30930
rect 26100 30090 26220 30210
rect 28620 31410 28740 31530
rect 27660 30270 27780 30390
rect 28140 31110 28260 31230
rect 40860 31410 40980 31530
rect 29700 31050 29820 31170
rect 29580 30810 29700 30930
rect 30900 30990 31020 31110
rect 31200 30990 31320 31110
rect 31620 31170 31740 31290
rect 31680 30930 31800 31050
rect 33180 31110 33300 31230
rect 32100 30990 32220 31110
rect 31890 30690 32010 30810
rect 29220 30090 29340 30210
rect 34620 31110 34740 31230
rect 33660 30270 33780 30390
rect 35100 30270 35220 30390
rect 36660 31050 36780 31170
rect 37740 31110 37860 31230
rect 36540 30810 36660 30930
rect 36180 30090 36300 30210
rect 39060 31050 39180 31170
rect 39180 30810 39300 30930
rect 38220 30270 38340 30390
rect 39540 30090 39660 30210
rect 41580 30270 41700 30390
rect 42060 31110 42180 31230
rect 43620 31050 43740 31170
rect 43500 30810 43620 30930
rect 44580 31050 44700 31170
rect 44700 30810 44820 30930
rect 43140 30090 43260 30210
rect 46140 30270 46260 30390
rect 45060 30090 45180 30210
rect 46620 31110 46740 31230
rect 48180 30990 48300 31110
rect 48660 31170 48780 31290
rect 48600 30930 48720 31050
rect 49080 30990 49200 31110
rect 49380 30990 49500 31110
rect 48390 30690 48510 30810
rect 7350 27390 7470 27510
rect 7140 27090 7260 27210
rect 7560 27150 7680 27270
rect 7620 26910 7740 27030
rect 8040 27090 8160 27210
rect 8340 27090 8460 27210
rect 8700 26970 8820 27090
rect 9180 27810 9300 27930
rect 11700 27990 11820 28110
rect 10230 27510 10350 27630
rect 9540 27090 9660 27210
rect 9840 27090 9960 27210
rect 10560 27330 10680 27450
rect 10260 26910 10380 27030
rect 10740 27090 10860 27210
rect 11340 27270 11460 27390
rect 11220 27030 11340 27150
rect 12060 26970 12180 27090
rect 12540 27810 12660 27930
rect 12780 26970 12900 27090
rect 13260 27810 13380 27930
rect 14130 27570 14250 27690
rect 13920 26970 14040 27090
rect 14460 27210 14580 27330
rect 15420 26970 15540 27090
rect 15900 27810 16020 27930
rect 16620 27810 16740 27930
rect 17100 26970 17220 27090
rect 18060 26970 18180 27090
rect 19380 27990 19500 28110
rect 18540 27810 18660 27930
rect 19740 27270 19860 27390
rect 19860 27030 19980 27150
rect 20940 26970 21060 27090
rect 21420 27810 21540 27930
rect 22140 26970 22260 27090
rect 22620 27810 22740 27930
rect 23580 26970 23700 27090
rect 24060 27810 24180 27930
rect 25020 26970 25140 27090
rect 25500 27810 25620 27930
rect 26460 26970 26580 27090
rect 28500 27990 28620 28110
rect 26940 27810 27060 27930
rect 30300 27810 30420 27930
rect 28860 27270 28980 27390
rect 28980 27030 29100 27150
rect 31860 27990 31980 28110
rect 30780 26970 30900 27090
rect 32220 27270 32340 27390
rect 32340 27030 32460 27150
rect 33270 27390 33390 27510
rect 33060 27090 33180 27210
rect 33480 27150 33600 27270
rect 33540 26910 33660 27030
rect 33960 27090 34080 27210
rect 34260 27090 34380 27210
rect 34860 26970 34980 27090
rect 35340 27810 35460 27930
rect 36060 26970 36180 27090
rect 36540 27810 36660 27930
rect 37500 27810 37620 27930
rect 37980 26970 38100 27090
rect 38700 26970 38820 27090
rect 39180 27810 39300 27930
rect 39990 27390 40110 27510
rect 39780 27090 39900 27210
rect 40200 27150 40320 27270
rect 40260 26910 40380 27030
rect 40680 27090 40800 27210
rect 40980 27090 41100 27210
rect 41580 26970 41700 27090
rect 43140 27990 43260 28110
rect 42060 27810 42180 27930
rect 45060 27990 45180 28110
rect 43500 27270 43620 27390
rect 43620 27030 43740 27150
rect 44700 27270 44820 27390
rect 44580 27030 44700 27150
rect 46500 27990 46620 28110
rect 46140 27270 46260 27390
rect 46020 27030 46140 27150
rect 47340 27510 47460 27630
rect 47610 27270 47730 27390
rect 48180 27450 48300 27570
rect 48060 27210 48180 27330
rect 48540 26970 48660 27090
rect 49020 27810 49140 27930
rect 49860 27990 49980 28110
rect 49500 27270 49620 27390
rect 49380 27030 49500 27150
rect 46860 26670 46980 26790
rect 12090 25410 12210 25530
rect 5460 24990 5580 25110
rect 5940 25170 6060 25290
rect 7020 25110 7140 25230
rect 5880 24930 6000 25050
rect 6360 24990 6480 25110
rect 6660 24990 6780 25110
rect 5670 24690 5790 24810
rect 7500 24270 7620 24390
rect 8340 25050 8460 25170
rect 8700 25110 8820 25230
rect 8220 24810 8340 24930
rect 7860 24090 7980 24210
rect 9540 24990 9660 25110
rect 10020 25170 10140 25290
rect 9960 24930 10080 25050
rect 10440 24990 10560 25110
rect 10740 24990 10860 25110
rect 9750 24690 9870 24810
rect 13980 25410 14100 25530
rect 12540 24870 12660 24990
rect 12660 24630 12780 24750
rect 9180 24270 9300 24390
rect 30540 25410 30660 25530
rect 15540 25050 15660 25170
rect 15420 24810 15540 24930
rect 15060 24090 15180 24210
rect 20700 24270 20820 24390
rect 21180 25110 21300 25230
rect 23100 25110 23220 25230
rect 25620 24990 25740 25110
rect 25920 24990 26040 25110
rect 26340 25170 26460 25290
rect 26400 24930 26520 25050
rect 26820 24990 26940 25110
rect 26610 24690 26730 24810
rect 23580 24270 23700 24390
rect 28500 25050 28620 25170
rect 28380 24810 28500 24930
rect 28020 24090 28140 24210
rect 32460 25410 32580 25530
rect 31620 25050 31740 25170
rect 31500 24810 31620 24930
rect 31140 24090 31260 24210
rect 43260 25410 43380 25530
rect 33180 25110 33300 25230
rect 34620 25110 34740 25230
rect 33660 24270 33780 24390
rect 36060 25110 36180 25230
rect 35100 24270 35220 24390
rect 37500 25110 37620 25230
rect 36540 24270 36660 24390
rect 38940 25110 39060 25230
rect 37980 24270 38100 24390
rect 40380 25110 40500 25230
rect 39420 24270 39540 24390
rect 41820 25110 41940 25230
rect 40860 24270 40980 24390
rect 44460 25410 44580 25530
rect 43740 24570 43860 24690
rect 42300 24270 42420 24390
rect 47940 24990 48060 25110
rect 48420 25170 48540 25290
rect 48360 24930 48480 25050
rect 48840 24990 48960 25110
rect 49140 24990 49260 25110
rect 48150 24690 48270 24810
rect 5670 21390 5790 21510
rect 5460 21090 5580 21210
rect 5880 21150 6000 21270
rect 5940 20910 6060 21030
rect 6360 21090 6480 21210
rect 6660 21090 6780 21210
rect 8220 20970 8340 21090
rect 8700 21810 8820 21930
rect 9660 20970 9780 21090
rect 11220 21990 11340 22110
rect 10140 21810 10260 21930
rect 11580 21270 11700 21390
rect 11700 21030 11820 21150
rect 14550 21390 14670 21510
rect 14340 21090 14460 21210
rect 14760 21150 14880 21270
rect 14820 20910 14940 21030
rect 15240 21090 15360 21210
rect 15540 21090 15660 21210
rect 18060 20970 18180 21090
rect 18540 21810 18660 21930
rect 22260 21990 22380 22110
rect 19890 21390 20010 21510
rect 18900 21090 19020 21210
rect 19200 21090 19320 21210
rect 19680 21150 19800 21270
rect 19620 20910 19740 21030
rect 21570 21390 21690 21510
rect 20100 21090 20220 21210
rect 20580 21090 20700 21210
rect 20880 21090 21000 21210
rect 21360 21150 21480 21270
rect 21300 20910 21420 21030
rect 21780 21090 21900 21210
rect 22620 21270 22740 21390
rect 22740 21030 22860 21150
rect 17100 20670 17220 20790
rect 26340 21990 26460 22110
rect 28020 21990 28140 22110
rect 26700 21270 26820 21390
rect 26820 21030 26940 21150
rect 28380 21270 28500 21390
rect 28500 21030 28620 21150
rect 29100 20970 29220 21090
rect 29580 21810 29700 21930
rect 30900 21990 31020 22110
rect 30540 21270 30660 21390
rect 30420 21030 30540 21150
rect 31980 20970 32100 21090
rect 32460 21810 32580 21930
rect 33180 20970 33300 21090
rect 33660 21810 33780 21930
rect 34620 20970 34740 21090
rect 35100 21810 35220 21930
rect 35820 20970 35940 21090
rect 36300 21810 36420 21930
rect 39060 21990 39180 22110
rect 37110 21390 37230 21510
rect 36900 21090 37020 21210
rect 37320 21150 37440 21270
rect 37380 20910 37500 21030
rect 37800 21090 37920 21210
rect 38100 21090 38220 21210
rect 39420 21270 39540 21390
rect 39540 21030 39660 21150
rect 40380 20970 40500 21090
rect 41700 21990 41820 22110
rect 40860 21810 40980 21930
rect 42060 21270 42180 21390
rect 42180 21030 42300 21150
rect 25020 20670 25140 20790
rect 43260 20670 43380 20790
rect 43740 21510 43860 21630
rect 44550 21390 44670 21510
rect 44340 21090 44460 21210
rect 44760 21150 44880 21270
rect 47010 21390 47130 21510
rect 44820 20910 44940 21030
rect 45240 21090 45360 21210
rect 45540 21090 45660 21210
rect 46020 21090 46140 21210
rect 46320 21090 46440 21210
rect 46800 21150 46920 21270
rect 46740 20910 46860 21030
rect 47220 21090 47340 21210
rect 48780 21510 48900 21630
rect 49050 21270 49170 21390
rect 49620 21450 49740 21570
rect 49500 21210 49620 21330
rect 47580 20670 47700 20790
rect 6180 19050 6300 19170
rect 6060 18810 6180 18930
rect 9060 18990 9180 19110
rect 9360 18990 9480 19110
rect 9780 19170 9900 19290
rect 9840 18930 9960 19050
rect 10260 18990 10380 19110
rect 11700 18990 11820 19110
rect 10050 18690 10170 18810
rect 12180 19170 12300 19290
rect 11880 18750 12000 18870
rect 12600 18990 12720 19110
rect 12900 18990 13020 19110
rect 13620 18990 13740 19110
rect 12210 18570 12330 18690
rect 14100 19170 14220 19290
rect 14040 18930 14160 19050
rect 14520 18990 14640 19110
rect 14820 18990 14940 19110
rect 13830 18690 13950 18810
rect 15660 18870 15780 18990
rect 15540 18630 15660 18750
rect 16110 19410 16230 19530
rect 27420 19410 27540 19530
rect 5700 18090 5820 18210
rect 18420 19050 18540 19170
rect 19500 19110 19620 19230
rect 18300 18810 18420 18930
rect 17940 18090 18060 18210
rect 20940 19110 21060 19230
rect 19980 18270 20100 18390
rect 22140 19110 22260 19230
rect 21420 18270 21540 18390
rect 23580 19110 23700 19230
rect 22620 18270 22740 18390
rect 24660 18990 24780 19110
rect 25140 19170 25260 19290
rect 25080 18930 25200 19050
rect 25560 18990 25680 19110
rect 25860 18990 25980 19110
rect 24870 18690 24990 18810
rect 26340 19050 26460 19170
rect 26460 18810 26580 18930
rect 24060 18270 24180 18390
rect 26820 18090 26940 18210
rect 36810 19410 36930 19530
rect 28980 19050 29100 19170
rect 30540 19110 30660 19230
rect 28860 18810 28980 18930
rect 28500 18090 28620 18210
rect 31980 19110 32100 19230
rect 31020 18270 31140 18390
rect 33300 19050 33420 19170
rect 33420 18810 33540 18930
rect 32460 18270 32580 18390
rect 35820 19110 35940 19230
rect 33780 18090 33900 18210
rect 41580 19410 41700 19530
rect 37260 18870 37380 18990
rect 37380 18630 37500 18750
rect 37980 19110 38100 19230
rect 36300 18270 36420 18390
rect 38940 19110 39060 19230
rect 38460 18270 38580 18390
rect 40380 19110 40500 19230
rect 39420 18270 39540 18390
rect 40860 18270 40980 18390
rect 47580 19410 47700 19530
rect 43020 18870 43140 18990
rect 42900 18630 43020 18750
rect 43470 18810 43590 18930
rect 44580 19050 44700 19170
rect 44700 18810 44820 18930
rect 43740 18570 43860 18690
rect 46140 19110 46260 19230
rect 45060 18090 45180 18210
rect 49140 19050 49260 19170
rect 49260 18810 49380 18930
rect 48060 18570 48180 18690
rect 46620 18270 46740 18390
rect 49620 18090 49740 18210
rect 6300 14970 6420 15090
rect 6780 15810 6900 15930
rect 8070 15390 8190 15510
rect 7860 15090 7980 15210
rect 8280 15150 8400 15270
rect 9750 15390 9870 15510
rect 8340 14910 8460 15030
rect 8760 15090 8880 15210
rect 9060 15090 9180 15210
rect 9540 15090 9660 15210
rect 9960 15150 10080 15270
rect 11730 15510 11850 15630
rect 11400 15330 11520 15450
rect 10020 14910 10140 15030
rect 10440 15090 10560 15210
rect 10740 15090 10860 15210
rect 11220 15090 11340 15210
rect 13890 15510 14010 15630
rect 13560 15330 13680 15450
rect 11700 14910 11820 15030
rect 12120 15090 12240 15210
rect 12420 15090 12540 15210
rect 13380 15090 13500 15210
rect 15270 15390 15390 15510
rect 13860 14910 13980 15030
rect 14280 15090 14400 15210
rect 14580 15090 14700 15210
rect 15060 15090 15180 15210
rect 15480 15150 15600 15270
rect 15540 14910 15660 15030
rect 15960 15090 16080 15210
rect 16260 15090 16380 15210
rect 16740 15450 16860 15570
rect 16860 15210 16980 15330
rect 18180 15990 18300 16110
rect 18540 15270 18660 15390
rect 18660 15030 18780 15150
rect 19260 14970 19380 15090
rect 19740 15810 19860 15930
rect 21300 15990 21420 16110
rect 22260 15990 22380 16110
rect 20940 15270 21060 15390
rect 20820 15030 20940 15150
rect 22620 15270 22740 15390
rect 22740 15030 22860 15150
rect 23580 14970 23700 15090
rect 24060 15810 24180 15930
rect 24780 15810 24900 15930
rect 26850 15390 26970 15510
rect 25860 15090 25980 15210
rect 26160 15090 26280 15210
rect 26640 15150 26760 15270
rect 25260 14970 25380 15090
rect 26580 14910 26700 15030
rect 27060 15090 27180 15210
rect 27900 14970 28020 15090
rect 28380 15810 28500 15930
rect 29100 14970 29220 15090
rect 29580 15810 29700 15930
rect 32220 15810 32340 15930
rect 31410 15390 31530 15510
rect 30420 15090 30540 15210
rect 30720 15090 30840 15210
rect 31200 15150 31320 15270
rect 31140 14910 31260 15030
rect 31620 15090 31740 15210
rect 32700 14970 32820 15090
rect 33180 14970 33300 15090
rect 33660 15810 33780 15930
rect 34620 14970 34740 15090
rect 35100 15810 35220 15930
rect 36660 15990 36780 16110
rect 36300 15270 36420 15390
rect 36180 15030 36300 15150
rect 37740 14970 37860 15090
rect 38220 15810 38340 15930
rect 45060 15990 45180 16110
rect 39810 15390 39930 15510
rect 38820 15090 38940 15210
rect 39120 15090 39240 15210
rect 39600 15150 39720 15270
rect 39540 14910 39660 15030
rect 41910 15390 42030 15510
rect 40020 15090 40140 15210
rect 41700 15090 41820 15210
rect 42120 15150 42240 15270
rect 42180 14910 42300 15030
rect 42600 15090 42720 15210
rect 42900 15090 43020 15210
rect 44700 15270 44820 15390
rect 44580 15030 44700 15150
rect 46140 14970 46260 15090
rect 46620 15810 46740 15930
rect 47580 15810 47700 15930
rect 49620 15990 49740 16110
rect 49260 15270 49380 15390
rect 48060 14970 48180 15090
rect 49140 15030 49260 15150
rect 17310 14670 17430 14790
rect 17820 14670 17940 14790
rect 6780 12270 6900 12390
rect 7260 13110 7380 13230
rect 9060 13050 9180 13170
rect 9180 12810 9300 12930
rect 10860 13110 10980 13230
rect 9660 12810 9780 12930
rect 9900 12870 10020 12990
rect 11340 12270 11460 12390
rect 12660 13050 12780 13170
rect 15900 13110 16020 13230
rect 12540 12810 12660 12930
rect 12180 12090 12300 12210
rect 16380 12270 16500 12390
rect 17220 13050 17340 13170
rect 17100 12810 17220 12930
rect 17700 12990 17820 13110
rect 18180 13170 18300 13290
rect 18120 12930 18240 13050
rect 18600 12990 18720 13110
rect 18900 12990 19020 13110
rect 19380 12990 19500 13110
rect 19680 12990 19800 13110
rect 20100 13170 20220 13290
rect 17910 12690 18030 12810
rect 20580 12990 20700 13110
rect 20400 12750 20520 12870
rect 20070 12570 20190 12690
rect 22020 12990 22140 13110
rect 22500 13170 22620 13290
rect 22200 12750 22320 12870
rect 22920 12990 23040 13110
rect 23220 12990 23340 13110
rect 22530 12570 22650 12690
rect 25140 13050 25260 13170
rect 25260 12810 25380 12930
rect 16740 12090 16860 12210
rect 26700 13110 26820 13230
rect 25620 12090 25740 12210
rect 29220 13050 29340 13170
rect 29340 12810 29460 12930
rect 27180 12270 27300 12390
rect 30900 13050 31020 13170
rect 30780 12810 30900 12930
rect 29700 12090 29820 12210
rect 30420 12090 30540 12210
rect 31980 12270 32100 12390
rect 32460 13110 32580 13230
rect 33060 12990 33180 13110
rect 33540 13170 33660 13290
rect 33480 12930 33600 13050
rect 33960 12990 34080 13110
rect 34260 12990 34380 13110
rect 33270 12690 33390 12810
rect 34740 13050 34860 13170
rect 34860 12810 34980 12930
rect 36060 13110 36180 13230
rect 35220 12090 35340 12210
rect 37500 13110 37620 13230
rect 36540 12270 36660 12390
rect 38940 13110 39060 13230
rect 37980 12270 38100 12390
rect 39420 12270 39540 12390
rect 40740 13050 40860 13170
rect 40620 12810 40740 12930
rect 41580 12870 41700 12990
rect 42120 13110 42240 13230
rect 43260 13110 43380 13230
rect 40260 12090 40380 12210
rect 41910 12510 42030 12630
rect 44580 13050 44700 13170
rect 44700 12810 44820 12930
rect 43740 12270 43860 12390
rect 46140 13110 46260 13230
rect 45060 12090 45180 12210
rect 47700 13050 47820 13170
rect 47820 12810 47940 12930
rect 46620 12270 46740 12390
rect 49260 12270 49380 12390
rect 48180 12090 48300 12210
rect 49740 13110 49860 13230
rect 5700 9990 5820 10110
rect 6060 9270 6180 9390
rect 6180 9030 6300 9150
rect 6780 8970 6900 9090
rect 7260 9810 7380 9930
rect 8070 9390 8190 9510
rect 7860 9090 7980 9210
rect 8280 9150 8400 9270
rect 8340 8910 8460 9030
rect 8760 9090 8880 9210
rect 9060 9090 9180 9210
rect 10050 9570 10170 9690
rect 11340 9810 11460 9930
rect 9840 8970 9960 9090
rect 10380 9210 10500 9330
rect 14070 9390 14190 9510
rect 13860 9090 13980 9210
rect 11820 8970 11940 9090
rect 14280 9150 14400 9270
rect 14340 8910 14460 9030
rect 14760 9090 14880 9210
rect 15060 9090 15180 9210
rect 16380 8970 16500 9090
rect 16860 9810 16980 9930
rect 21180 9810 21300 9930
rect 17970 9510 18090 9630
rect 17640 9330 17760 9450
rect 17460 9090 17580 9210
rect 20370 9390 20490 9510
rect 17940 8910 18060 9030
rect 18360 9090 18480 9210
rect 18660 9090 18780 9210
rect 19380 9090 19500 9210
rect 19680 9090 19800 9210
rect 20160 9150 20280 9270
rect 20100 8910 20220 9030
rect 20580 9090 20700 9210
rect 23010 9390 23130 9510
rect 22020 9090 22140 9210
rect 22320 9090 22440 9210
rect 22800 9150 22920 9270
rect 21660 8970 21780 9090
rect 22740 8910 22860 9030
rect 23220 9090 23340 9210
rect 23820 8970 23940 9090
rect 24300 9810 24420 9930
rect 25830 9390 25950 9510
rect 25620 9090 25740 9210
rect 26040 9150 26160 9270
rect 26100 8910 26220 9030
rect 26520 9090 26640 9210
rect 26820 9090 26940 9210
rect 27900 8970 28020 9090
rect 28380 9810 28500 9930
rect 32340 9990 32460 10110
rect 31980 9270 32100 9390
rect 31860 9030 31980 9150
rect 33990 9510 34110 9630
rect 33300 9090 33420 9210
rect 33600 9090 33720 9210
rect 34320 9330 34440 9450
rect 34020 8910 34140 9030
rect 34500 9090 34620 9210
rect 35970 9570 36090 9690
rect 35760 8970 35880 9090
rect 29580 8670 29700 8790
rect 30540 8670 30660 8790
rect 36300 9210 36420 9330
rect 36780 8970 36900 9090
rect 37260 9810 37380 9930
rect 38130 9570 38250 9690
rect 39540 9990 39660 10110
rect 37920 8970 38040 9090
rect 38460 9210 38580 9330
rect 39180 9270 39300 9390
rect 39060 9030 39180 9150
rect 40380 8970 40500 9090
rect 40860 9810 40980 9930
rect 41580 8970 41700 9090
rect 42060 9810 42180 9930
rect 47580 9810 47700 9930
rect 42870 9390 42990 9510
rect 42660 9090 42780 9210
rect 43080 9150 43200 9270
rect 45510 9390 45630 9510
rect 43140 8910 43260 9030
rect 43560 9090 43680 9210
rect 43860 9090 43980 9210
rect 45300 9090 45420 9210
rect 45720 9150 45840 9270
rect 45780 8910 45900 9030
rect 46200 9090 46320 9210
rect 46500 9090 46620 9210
rect 49020 9810 49140 9930
rect 48060 8970 48180 9090
rect 49500 8970 49620 9090
rect 8220 7410 8340 7530
rect 5700 6990 5820 7110
rect 6000 6990 6120 7110
rect 6420 7170 6540 7290
rect 6480 6930 6600 7050
rect 6900 6990 7020 7110
rect 6690 6690 6810 6810
rect 9300 7050 9420 7170
rect 9900 7110 10020 7230
rect 9180 6810 9300 6930
rect 8820 6090 8940 6210
rect 10380 6270 10500 6390
rect 11460 7050 11580 7170
rect 12300 7110 12420 7230
rect 11340 6810 11460 6930
rect 10980 6090 11100 6210
rect 13980 6870 14100 6990
rect 13860 6630 13980 6750
rect 14430 7410 14550 7530
rect 15420 7410 15540 7530
rect 18060 7410 18180 7530
rect 15900 6570 16020 6690
rect 43260 7410 43380 7530
rect 20700 7110 20820 7230
rect 18540 6570 18660 6690
rect 12780 6270 12900 6390
rect 23340 7110 23460 7230
rect 21180 6270 21300 6390
rect 25860 6990 25980 7110
rect 26340 7170 26460 7290
rect 27900 7110 28020 7230
rect 26040 6750 26160 6870
rect 26760 6990 26880 7110
rect 27060 6990 27180 7110
rect 26370 6570 26490 6690
rect 23820 6270 23940 6390
rect 29100 7110 29220 7230
rect 28380 6270 28500 6390
rect 30180 6990 30300 7110
rect 30660 7170 30780 7290
rect 30600 6930 30720 7050
rect 31080 6990 31200 7110
rect 31380 6990 31500 7110
rect 30390 6690 30510 6810
rect 32100 7050 32220 7170
rect 32220 6810 32340 6930
rect 29580 6270 29700 6390
rect 33180 7110 33300 7230
rect 32580 6090 32700 6210
rect 33660 6270 33780 6390
rect 34620 6270 34740 6390
rect 35100 7110 35220 7230
rect 36060 7110 36180 7230
rect 36540 6270 36660 6390
rect 38100 7050 38220 7170
rect 38940 7110 39060 7230
rect 37980 6810 38100 6930
rect 37620 6090 37740 6210
rect 40380 7110 40500 7230
rect 39420 6270 39540 6390
rect 46620 7410 46740 7530
rect 44700 6870 44820 6990
rect 43740 6570 43860 6690
rect 44580 6630 44700 6750
rect 45150 6810 45270 6930
rect 45420 6570 45540 6690
rect 40860 6270 40980 6390
rect 47940 7050 48060 7170
rect 47820 6810 47940 6930
rect 47460 6090 47580 6210
<< metal1 >>
rect 1155 48076 54240 48135
rect 1155 47204 1214 48076
rect 2086 47204 53310 48076
rect 54180 47204 54240 48076
rect 1155 47145 54240 47204
rect 15180 46590 15300 46710
rect 15420 46605 32940 46695
rect 3135 46096 52260 46155
rect 3135 45224 3194 46096
rect 4066 45224 51330 46096
rect 52200 45224 52260 46096
rect 3135 45165 52260 45224
rect 3135 44160 52260 44190
rect 3135 44040 3194 44160
rect 4066 44040 5220 44160
rect 5340 44040 5460 44160
rect 5580 44040 5940 44160
rect 6060 44040 6420 44160
rect 6540 44040 6660 44160
rect 6780 44040 7140 44160
rect 7260 44040 7380 44160
rect 7500 44040 7620 44160
rect 7740 44040 8100 44160
rect 8220 44040 8580 44160
rect 8700 44040 8820 44160
rect 8940 44040 9300 44160
rect 9420 44040 9780 44160
rect 9900 44040 10260 44160
rect 10380 44040 10500 44160
rect 10620 44040 10740 44160
rect 10860 44040 10980 44160
rect 11100 44040 11460 44160
rect 11580 44040 11700 44160
rect 11820 44040 11940 44160
rect 12060 44040 12180 44160
rect 12300 44040 12420 44160
rect 12540 44040 12900 44160
rect 13020 44040 13140 44160
rect 13260 44040 13380 44160
rect 13500 44040 13620 44160
rect 13740 44040 14100 44160
rect 14220 44040 14580 44160
rect 14700 44040 14820 44160
rect 14940 44040 15060 44160
rect 15180 44040 15300 44160
rect 15420 44040 15780 44160
rect 15900 44040 16020 44160
rect 16140 44040 16260 44160
rect 16380 44040 16500 44160
rect 16620 44040 16740 44160
rect 16860 44040 16980 44160
rect 17100 44040 17460 44160
rect 17580 44040 17940 44160
rect 18060 44040 18180 44160
rect 18300 44040 18420 44160
rect 18540 44040 18660 44160
rect 18780 44040 18900 44160
rect 19020 44040 19140 44160
rect 19260 44040 19380 44160
rect 19500 44040 19860 44160
rect 19980 44040 20340 44160
rect 20460 44040 20820 44160
rect 20940 44040 21060 44160
rect 21180 44040 21540 44160
rect 21660 44040 21780 44160
rect 21900 44040 22020 44160
rect 22140 44040 22260 44160
rect 22380 44040 22500 44160
rect 22620 44040 22980 44160
rect 23100 44040 23460 44160
rect 23580 44040 23940 44160
rect 24060 44040 24180 44160
rect 24300 44040 24420 44160
rect 24540 44040 24660 44160
rect 24780 44040 24900 44160
rect 25020 44040 25380 44160
rect 25500 44040 25860 44160
rect 25980 44040 26100 44160
rect 26220 44040 26340 44160
rect 26460 44040 26580 44160
rect 26700 44040 27060 44160
rect 27180 44040 27300 44160
rect 27420 44040 27540 44160
rect 27660 44040 27780 44160
rect 27900 44040 28260 44160
rect 28380 44040 28740 44160
rect 28860 44040 28980 44160
rect 29100 44040 29460 44160
rect 29580 44040 29700 44160
rect 29820 44040 29940 44160
rect 30060 44040 30180 44160
rect 30300 44040 30660 44160
rect 30780 44040 31140 44160
rect 31260 44040 31380 44160
rect 31500 44040 31620 44160
rect 31740 44040 32100 44160
rect 32220 44040 32580 44160
rect 32700 44040 32820 44160
rect 32940 44040 33060 44160
rect 33180 44040 33300 44160
rect 33420 44040 33780 44160
rect 33900 44040 34020 44160
rect 34140 44040 34260 44160
rect 34380 44040 34500 44160
rect 34620 44040 34980 44160
rect 35100 44040 35220 44160
rect 35340 44040 35460 44160
rect 35580 44040 35700 44160
rect 35820 44040 36180 44160
rect 36300 44040 36660 44160
rect 36780 44040 37140 44160
rect 37260 44040 37380 44160
rect 37500 44040 37620 44160
rect 37740 44040 38100 44160
rect 38220 44040 38580 44160
rect 38700 44040 38820 44160
rect 38940 44040 39060 44160
rect 39180 44040 39300 44160
rect 39420 44040 39540 44160
rect 39660 44040 40020 44160
rect 40140 44040 40500 44160
rect 40620 44040 40980 44160
rect 41100 44040 41220 44160
rect 41340 44040 41460 44160
rect 41580 44040 41700 44160
rect 41820 44040 42180 44160
rect 42300 44040 42420 44160
rect 42540 44040 42660 44160
rect 42780 44040 42900 44160
rect 43020 44040 43380 44160
rect 43500 44040 43860 44160
rect 43980 44040 44100 44160
rect 44220 44040 44580 44160
rect 44700 44040 45540 44160
rect 45660 44040 46020 44160
rect 46140 44040 46500 44160
rect 46620 44040 46980 44160
rect 47100 44040 47220 44160
rect 47340 44040 47700 44160
rect 47820 44040 48180 44160
rect 48300 44040 48660 44160
rect 48780 44040 48900 44160
rect 49020 44040 49140 44160
rect 49260 44040 49380 44160
rect 49500 44040 49620 44160
rect 49740 44040 49860 44160
rect 49980 44040 50100 44160
rect 50220 44040 51330 44160
rect 52200 44040 52260 44160
rect 3135 44010 52260 44040
rect 6060 43890 6180 44010
rect 6780 43920 6900 44010
rect 6060 43440 6180 43470
rect 5940 43320 6300 43350
rect 7020 43320 7170 43410
rect 7500 43695 7620 43710
rect 7500 43605 7740 43695
rect 7500 43590 7620 43605
rect 8220 43890 8340 44010
rect 9210 43920 9330 44010
rect 8220 43440 8340 43470
rect 8100 43320 8460 43350
rect 9180 43890 9330 43920
rect 9180 43410 9330 43440
rect 9600 43860 9840 43920
rect 9600 43440 9660 43860
rect 9780 43440 9840 43860
rect 9600 43380 9840 43440
rect 10110 43890 10260 44010
rect 10860 43920 10980 44010
rect 11340 43920 11460 44010
rect 10110 43410 10260 43440
rect 5610 43110 5700 43320
rect 5850 43260 6390 43320
rect 5580 43095 5970 43110
rect 5460 43005 5970 43095
rect 6300 43095 6420 43110
rect 6540 43095 6660 43110
rect 6300 43050 6660 43095
rect 6180 43020 6660 43050
rect 5580 42990 5970 43005
rect 6300 43005 6660 43020
rect 6300 42990 6420 43005
rect 6540 42990 6660 43005
rect 6780 42990 6900 43110
rect 5580 42480 5700 42510
rect 5880 42480 5970 42990
rect 6795 42810 6885 42990
rect 6060 42795 6180 42810
rect 6780 42795 6900 42810
rect 6060 42705 6900 42795
rect 6060 42690 6180 42705
rect 6780 42690 6900 42705
rect 6540 42495 6660 42510
rect 7020 42495 7140 43320
rect 7770 43110 7860 43320
rect 8010 43260 8550 43320
rect 8940 43230 9210 43320
rect 7740 42990 8130 43110
rect 8460 43095 8580 43110
rect 8460 43050 8940 43095
rect 8340 43020 8940 43050
rect 8460 43005 8940 43020
rect 8460 42990 8580 43005
rect 9750 43080 9840 43380
rect 12300 43920 12420 44010
rect 12780 43920 12900 44010
rect 10260 43230 10500 43320
rect 9180 43050 9270 43080
rect 5580 42390 5790 42480
rect 5880 42466 6030 42480
rect 5880 42390 5910 42466
rect 5700 42210 5790 42390
rect 5670 41866 5790 41880
rect 5670 41190 5790 41294
rect 5910 41280 6030 41294
rect 6300 42466 6420 42480
rect 6540 42405 7140 42495
rect 6540 42390 6660 42405
rect 6300 41190 6420 41294
rect 6780 41866 6900 41880
rect 6780 41190 6900 41294
rect 7020 41866 7140 42405
rect 7740 42480 7860 42510
rect 8040 42480 8130 42990
rect 9180 42960 9480 43050
rect 9690 42990 9840 43080
rect 9960 43110 10050 43170
rect 11100 43110 11190 43620
rect 11340 43395 11460 43410
rect 12300 43395 12420 43410
rect 11340 43305 12420 43395
rect 11340 43290 11460 43305
rect 12300 43290 12420 43305
rect 12540 43110 12630 43620
rect 13980 43890 14100 44010
rect 15420 43920 15540 44010
rect 13980 43440 14100 43470
rect 13860 43320 14220 43350
rect 15660 43320 15810 43410
rect 17340 43890 17460 44010
rect 17340 43440 17460 43470
rect 17220 43320 17580 43350
rect 19500 43890 19650 44010
rect 20430 43920 20550 44010
rect 21180 43920 21300 44010
rect 22890 43920 23010 44010
rect 19500 43410 19650 43440
rect 19920 43860 20160 43920
rect 19920 43440 19980 43860
rect 20100 43440 20160 43860
rect 19920 43380 20160 43440
rect 20430 43890 20580 43920
rect 20430 43410 20580 43440
rect 13770 43260 14310 43320
rect 10380 42990 10500 43110
rect 11100 43095 11220 43110
rect 10740 43005 11220 43095
rect 11100 42990 11220 43005
rect 11340 43095 11460 43110
rect 12540 43095 12660 43110
rect 11340 43005 12660 43095
rect 11340 42990 11460 43005
rect 12540 42990 12660 43005
rect 13740 43095 13860 43110
rect 12900 43050 13860 43095
rect 14460 43110 14550 43320
rect 12900 43020 13980 43050
rect 12900 43005 13860 43020
rect 13740 42990 13860 43005
rect 14190 42990 14220 43110
rect 14340 42990 14580 43110
rect 14700 43095 14820 43110
rect 15420 43095 15540 43110
rect 14700 43005 15540 43095
rect 14700 42990 14820 43005
rect 15420 42990 15540 43005
rect 9690 42810 9780 42990
rect 8220 42795 8340 42810
rect 8220 42705 8700 42795
rect 8220 42690 8340 42705
rect 9660 42690 9780 42810
rect 9690 42480 9780 42690
rect 11100 42480 11190 42990
rect 12300 42795 12420 42810
rect 11700 42705 12420 42795
rect 12300 42690 12420 42705
rect 12540 42480 12630 42990
rect 13980 42795 14100 42810
rect 13140 42705 14100 42795
rect 13980 42690 14100 42705
rect 14190 42480 14280 42990
rect 14460 42495 14580 42510
rect 15660 42495 15780 43320
rect 17130 43260 17670 43320
rect 17820 43110 17910 43320
rect 19260 43230 19500 43320
rect 19710 43110 19800 43170
rect 17220 43020 17340 43050
rect 17550 42990 17580 43110
rect 17700 42990 17940 43110
rect 17340 42690 17460 42810
rect 14460 42480 15780 42495
rect 7740 42390 7950 42480
rect 8040 42466 8190 42480
rect 8040 42390 8070 42466
rect 7860 42210 7950 42390
rect 7020 41280 7140 41294
rect 7260 41866 7380 41880
rect 7260 41190 7380 41294
rect 7830 41866 7950 41880
rect 7830 41190 7950 41294
rect 8070 41280 8190 41294
rect 8460 42466 8580 42480
rect 8460 41190 8580 41294
rect 8940 42466 9210 42480
rect 9060 42390 9210 42466
rect 9600 42466 9840 42480
rect 8940 41280 9060 41294
rect 9180 42210 9330 42270
rect 9180 41340 9194 42210
rect 9316 41340 9330 42210
rect 9180 41280 9330 41340
rect 9600 41294 9660 42466
rect 9780 41294 9840 42466
rect 10260 42466 10500 42480
rect 10260 42390 10380 42466
rect 9600 41280 9840 41294
rect 10110 42210 10260 42270
rect 10110 41340 10124 42210
rect 10246 41340 10260 42210
rect 9210 41190 9330 41280
rect 10110 41190 10260 41340
rect 10380 41280 10500 41294
rect 11070 42360 11220 42480
rect 10950 41280 11070 41310
rect 11340 41190 11460 41310
rect 12510 42360 12660 42480
rect 12390 41280 12510 41310
rect 12780 41190 12900 41310
rect 13740 42466 13860 42480
rect 13740 41190 13860 41294
rect 14130 42466 14280 42480
rect 14250 42390 14280 42466
rect 14370 42405 15780 42480
rect 14370 42390 14580 42405
rect 14370 42210 14460 42390
rect 14130 41280 14250 41294
rect 14370 41866 14490 41880
rect 14370 41190 14490 41294
rect 15420 41866 15540 41880
rect 15420 41190 15540 41294
rect 15660 41866 15780 42405
rect 15900 42390 16020 42510
rect 17550 42480 17640 42990
rect 19920 42870 20010 43380
rect 21180 43620 21300 43650
rect 20340 43170 20400 43260
rect 20610 43230 20820 43320
rect 21180 43395 21300 43410
rect 21060 43305 21300 43395
rect 21180 43290 21300 43305
rect 20310 43110 20400 43170
rect 20310 43020 20580 43110
rect 20700 42990 20820 43110
rect 19860 42810 20010 42870
rect 19740 42795 20010 42810
rect 18180 42780 20010 42795
rect 20130 42870 20220 42960
rect 20130 42780 20400 42870
rect 18180 42705 19950 42780
rect 20700 42795 20820 42810
rect 21420 42795 21540 43650
rect 22860 43890 23010 43920
rect 22860 43410 23010 43440
rect 23280 43860 23520 43920
rect 23280 43440 23340 43860
rect 23460 43440 23520 43860
rect 23280 43380 23520 43440
rect 23790 43890 23940 44010
rect 23790 43410 23940 43440
rect 22620 43230 22890 43320
rect 23430 43080 23520 43380
rect 25500 43890 25620 44010
rect 26700 43920 26820 44010
rect 25500 43440 25620 43470
rect 25380 43320 25740 43350
rect 26940 43320 27090 43410
rect 28140 43890 28260 44010
rect 29100 43920 29220 44010
rect 28140 43440 28260 43470
rect 28020 43320 28380 43350
rect 29340 43320 29490 43410
rect 30540 43890 30660 44010
rect 30540 43440 30660 43470
rect 30420 43320 30780 43350
rect 31140 43605 31500 43695
rect 31980 43890 32100 44010
rect 33660 43920 33780 44010
rect 31980 43440 32100 43470
rect 31860 43320 32220 43350
rect 33390 43320 33540 43410
rect 34620 43920 34740 44010
rect 35100 43920 35220 44010
rect 36090 43920 36210 44010
rect 23940 43230 24180 43320
rect 22860 43050 22950 43080
rect 22860 42960 23160 43050
rect 23370 42990 23520 43080
rect 23640 43110 23730 43170
rect 25050 43110 25140 43320
rect 25290 43260 25830 43320
rect 24060 43095 24180 43110
rect 25020 43095 25410 43110
rect 24060 43005 25410 43095
rect 25620 43020 25740 43050
rect 24060 42990 24180 43005
rect 25020 42990 25410 43005
rect 26700 43095 26820 43110
rect 25995 43005 26820 43095
rect 23370 42810 23460 42990
rect 19740 42690 19950 42705
rect 20700 42705 21540 42795
rect 20700 42690 20820 42705
rect 17820 42495 17940 42510
rect 17820 42480 18780 42495
rect 17100 42466 17220 42480
rect 15660 41280 15780 41294
rect 15900 41866 16020 41880
rect 15900 41190 16020 41294
rect 17100 41190 17220 41294
rect 17490 42466 17640 42480
rect 17610 42390 17640 42466
rect 17730 42405 18780 42480
rect 17730 42390 17940 42405
rect 19860 42480 19950 42690
rect 20190 42570 20580 42660
rect 20490 42480 20580 42570
rect 19260 42466 19500 42480
rect 17730 42210 17820 42390
rect 17490 41280 17610 41294
rect 17730 41866 17850 41880
rect 17730 41190 17850 41294
rect 19380 42390 19500 42466
rect 19860 42466 20160 42480
rect 19860 42390 19980 42466
rect 19260 41280 19380 41294
rect 19500 42210 19650 42270
rect 19500 41340 19514 42210
rect 19636 41340 19650 42210
rect 19500 41190 19650 41340
rect 19920 41294 19980 42390
rect 20100 41294 20160 42466
rect 20610 42466 20820 42480
rect 20610 42390 20700 42466
rect 19920 41280 20160 41294
rect 20430 42210 20580 42270
rect 20430 41340 20444 42210
rect 20566 41340 20580 42210
rect 20430 41280 20580 41340
rect 21420 41880 21540 42705
rect 23340 42690 23460 42810
rect 23370 42480 23460 42690
rect 25020 42480 25140 42510
rect 25320 42480 25410 42990
rect 25500 42795 25620 42810
rect 25995 42795 26085 43005
rect 26700 42990 26820 43005
rect 25500 42705 26220 42795
rect 25500 42690 25620 42705
rect 25980 42495 26100 42510
rect 26940 42495 27060 43320
rect 27930 43260 28470 43320
rect 27300 43005 27900 43095
rect 28620 43110 28710 43320
rect 28020 43020 28140 43050
rect 28350 42990 28740 43110
rect 28860 43095 28980 43110
rect 29100 43095 29220 43110
rect 28860 43005 29220 43095
rect 28860 42990 28980 43005
rect 29100 42990 29220 43005
rect 20700 41280 20820 41294
rect 20430 41190 20550 41280
rect 21180 41190 21300 41310
rect 21420 41280 21540 41310
rect 22620 42466 22890 42480
rect 22740 42390 22890 42466
rect 23280 42466 23520 42480
rect 22620 41280 22740 41294
rect 22860 42210 23010 42270
rect 22860 41340 22874 42210
rect 22996 41340 23010 42210
rect 22860 41280 23010 41340
rect 23280 41294 23340 42466
rect 23460 41294 23520 42466
rect 23940 42466 24180 42480
rect 23940 42390 24060 42466
rect 23280 41280 23520 41294
rect 23790 42210 23940 42270
rect 23790 41340 23804 42210
rect 23926 41340 23940 42210
rect 22890 41190 23010 41280
rect 23790 41190 23940 41340
rect 25020 42390 25230 42480
rect 25320 42466 25470 42480
rect 25320 42390 25350 42466
rect 25140 42210 25230 42390
rect 24060 41280 24180 41294
rect 25110 41866 25230 41880
rect 25110 41190 25230 41294
rect 25350 41280 25470 41294
rect 25740 42466 25860 42480
rect 25980 42405 27060 42495
rect 25980 42390 26100 42405
rect 25740 41190 25860 41294
rect 26700 41866 26820 41880
rect 26700 41190 26820 41294
rect 26940 41866 27060 42405
rect 28350 42480 28440 42990
rect 28620 42495 28740 42510
rect 29340 42495 29460 43320
rect 30330 43260 30870 43320
rect 30300 43095 30420 43110
rect 29700 43050 30420 43095
rect 31020 43110 31110 43320
rect 31770 43260 32310 43320
rect 29700 43020 30540 43050
rect 29700 43005 30420 43020
rect 30300 42990 30420 43005
rect 30750 42990 31140 43110
rect 31740 43095 31860 43110
rect 31380 43050 31860 43095
rect 32460 43110 32550 43320
rect 31380 43020 31980 43050
rect 31380 43005 31860 43020
rect 31740 42990 31860 43005
rect 32190 42990 32580 43110
rect 30540 42690 30660 42810
rect 28620 42480 29460 42495
rect 27900 42466 28020 42480
rect 26940 41280 27060 41294
rect 27180 41866 27300 41880
rect 27180 41190 27300 41294
rect 27900 41190 28020 41294
rect 28290 42466 28440 42480
rect 28410 42390 28440 42466
rect 28530 42405 29460 42480
rect 28530 42390 28740 42405
rect 28530 42210 28620 42390
rect 28290 41280 28410 41294
rect 28530 41866 28650 41880
rect 28530 41190 28650 41294
rect 29100 41866 29220 41880
rect 29100 41190 29220 41294
rect 29340 41866 29460 42405
rect 29580 42390 29700 42510
rect 30750 42480 30840 42990
rect 31980 42690 32100 42810
rect 31020 42495 31140 42510
rect 31500 42495 31620 42510
rect 31020 42480 31620 42495
rect 32190 42480 32280 42990
rect 33420 42795 33540 43320
rect 34890 43110 34980 43620
rect 36060 43890 36210 43920
rect 36060 43410 36210 43440
rect 36480 43860 36720 43920
rect 36480 43440 36540 43860
rect 36660 43440 36720 43860
rect 36480 43380 36720 43440
rect 36990 43890 37140 44010
rect 36990 43410 37140 43440
rect 35820 43230 36090 43320
rect 34860 43095 34980 43110
rect 34860 43005 35820 43095
rect 34860 42990 34980 43005
rect 36630 43080 36720 43380
rect 38220 43890 38340 44010
rect 38220 43440 38340 43470
rect 38100 43320 38460 43350
rect 39660 43890 39810 44010
rect 40590 43920 40710 44010
rect 41820 43920 41940 44010
rect 39660 43410 39810 43440
rect 40080 43860 40320 43920
rect 40080 43440 40140 43860
rect 40260 43440 40320 43860
rect 40080 43380 40320 43440
rect 40590 43890 40740 43920
rect 40590 43410 40740 43440
rect 37140 43230 37380 43320
rect 36060 43050 36150 43080
rect 32955 42705 33540 42795
rect 32460 42495 32580 42510
rect 32955 42495 33045 42705
rect 32460 42480 33045 42495
rect 30300 42466 30420 42480
rect 29340 41280 29460 41294
rect 29580 41866 29700 41880
rect 29580 41190 29700 41294
rect 30300 41190 30420 41294
rect 30690 42466 30840 42480
rect 30810 42390 30840 42466
rect 30930 42405 31620 42480
rect 30930 42390 31140 42405
rect 31500 42390 31620 42405
rect 31740 42466 31860 42480
rect 30930 42210 31020 42390
rect 30690 41280 30810 41294
rect 30930 41866 31050 41880
rect 30930 41190 31050 41294
rect 31740 41190 31860 41294
rect 32130 42466 32280 42480
rect 32250 42390 32280 42466
rect 32370 42405 33045 42480
rect 32370 42390 32580 42405
rect 32370 42210 32460 42390
rect 32130 41280 32250 41294
rect 32370 41866 32490 41880
rect 32370 41190 32490 41294
rect 33180 41866 33300 41880
rect 33180 41190 33300 41294
rect 33420 41866 33540 42705
rect 34890 42480 34980 42990
rect 36060 42960 36360 43050
rect 36570 42990 36720 43080
rect 36840 43110 36930 43170
rect 37770 43110 37860 43320
rect 38010 43260 38550 43320
rect 39420 43230 39660 43320
rect 37260 43095 37380 43110
rect 37740 43095 38130 43110
rect 37260 43005 38130 43095
rect 39870 43110 39960 43170
rect 38460 43050 38580 43110
rect 38340 43020 38580 43050
rect 37260 42990 37380 43005
rect 37740 42990 38130 43005
rect 38460 42990 38580 43020
rect 40080 43080 40170 43380
rect 41820 43620 41940 43650
rect 40710 43230 40980 43320
rect 41340 43395 41460 43410
rect 41820 43395 41940 43410
rect 41340 43305 41940 43395
rect 41340 43290 41460 43305
rect 41820 43290 41940 43305
rect 40080 42990 40230 43080
rect 40650 43050 40740 43080
rect 36570 42810 36660 42990
rect 35100 42795 35220 42810
rect 35100 42705 35340 42795
rect 35100 42690 35220 42705
rect 36540 42690 36660 42810
rect 36570 42480 36660 42690
rect 33420 41280 33540 41294
rect 33660 41866 33780 41880
rect 33660 41190 33780 41294
rect 34860 42360 35010 42480
rect 34620 41190 34740 41310
rect 35010 41280 35130 41310
rect 35820 42466 36090 42480
rect 35940 42390 36090 42466
rect 36480 42466 36720 42480
rect 35820 41280 35940 41294
rect 36060 42210 36210 42270
rect 36060 41340 36074 42210
rect 36196 41340 36210 42210
rect 36060 41280 36210 41340
rect 36480 41294 36540 42466
rect 36660 41294 36720 42466
rect 37140 42466 37380 42480
rect 37140 42390 37260 42466
rect 36480 41280 36720 41294
rect 36990 42210 37140 42270
rect 36990 41340 37004 42210
rect 37126 41340 37140 42210
rect 36090 41190 36210 41280
rect 36990 41190 37140 41340
rect 38040 42480 38130 42990
rect 40140 42810 40230 42990
rect 40440 42960 40740 43050
rect 40140 42690 40260 42810
rect 40140 42480 40230 42690
rect 42060 42795 42180 43650
rect 43260 43890 43380 44010
rect 43260 43440 43380 43470
rect 43140 43320 43500 43350
rect 44460 43890 44580 44010
rect 45420 43920 45540 44010
rect 45930 43920 46050 44010
rect 44460 43440 44580 43470
rect 44340 43320 44700 43350
rect 43050 43260 43590 43320
rect 43020 43095 43140 43110
rect 42420 43050 43140 43095
rect 43740 43110 43830 43320
rect 44250 43260 44790 43320
rect 42420 43020 43260 43050
rect 43470 43095 43860 43110
rect 44220 43095 44340 43110
rect 43470 43050 44340 43095
rect 44940 43110 45030 43320
rect 43470 43020 44460 43050
rect 42420 43005 43140 43020
rect 43020 42990 43140 43005
rect 43470 43005 44340 43020
rect 43470 42990 43860 43005
rect 44220 42990 44340 43005
rect 44670 42990 44940 43110
rect 43260 42795 43380 42810
rect 42060 42705 43380 42795
rect 37860 42210 37950 42480
rect 38040 42466 38190 42480
rect 38040 42390 38070 42466
rect 37260 41280 37380 41294
rect 37830 41866 37950 41880
rect 37830 41190 37950 41294
rect 38070 41280 38190 41294
rect 38460 42466 38580 42480
rect 38460 41190 38580 41294
rect 39420 42466 39660 42480
rect 39540 42390 39660 42466
rect 40080 42466 40320 42480
rect 39420 41280 39540 41294
rect 39660 42210 39810 42270
rect 39660 41340 39674 42210
rect 39796 41340 39810 42210
rect 39660 41190 39810 41340
rect 40080 41294 40140 42466
rect 40260 41294 40320 42466
rect 40710 42466 40980 42480
rect 40710 42390 40860 42466
rect 40080 41280 40320 41294
rect 40590 42210 40740 42270
rect 40590 41340 40604 42210
rect 40726 41340 40740 42210
rect 40590 41280 40740 41340
rect 42060 41880 42180 42705
rect 43260 42690 43380 42705
rect 43470 42480 43560 42990
rect 44460 42690 44580 42810
rect 43740 42495 43860 42510
rect 43740 42480 43980 42495
rect 40860 41280 40980 41294
rect 40590 41190 40710 41280
rect 41820 41190 41940 41310
rect 42060 41280 42180 41310
rect 43020 42466 43140 42480
rect 43020 41190 43140 41294
rect 43410 42466 43560 42480
rect 43530 42390 43560 42466
rect 43650 42405 43980 42480
rect 43650 42390 43860 42405
rect 44670 42480 44760 42990
rect 44940 42795 45060 42810
rect 45180 42795 45300 43650
rect 45420 43620 45540 43650
rect 45900 43890 46050 43920
rect 45900 43410 46050 43440
rect 46320 43860 46560 43920
rect 46320 43440 46380 43860
rect 46500 43440 46560 43860
rect 46320 43380 46560 43440
rect 46830 43890 46980 44010
rect 47610 43920 47730 44010
rect 46830 43410 46980 43440
rect 45660 43230 45930 43320
rect 45420 43095 45540 43110
rect 45660 43095 45780 43110
rect 45420 43005 45780 43095
rect 45420 42990 45540 43005
rect 45660 42990 45780 43005
rect 46470 43080 46560 43380
rect 46980 43230 47220 43320
rect 47580 43890 47730 43920
rect 47580 43410 47730 43440
rect 48000 43860 48240 43920
rect 48000 43440 48060 43860
rect 48180 43440 48240 43860
rect 48000 43380 48240 43440
rect 48510 43890 48660 44010
rect 48510 43410 48660 43440
rect 47340 43230 47610 43320
rect 45900 43050 45990 43080
rect 45900 42960 46200 43050
rect 46410 42990 46560 43080
rect 46680 43110 46770 43170
rect 48150 43080 48240 43380
rect 48660 43230 48900 43320
rect 47580 43050 47670 43080
rect 46410 42810 46500 42990
rect 47580 42960 47880 43050
rect 48090 42990 48240 43080
rect 48360 43110 48450 43170
rect 48090 42810 48180 42990
rect 44940 42705 45300 42795
rect 44940 42690 45060 42705
rect 44220 42466 44340 42480
rect 43650 42210 43740 42390
rect 43410 41280 43530 41294
rect 43650 41866 43770 41880
rect 43650 41190 43770 41294
rect 44220 41190 44340 41294
rect 44610 42466 44760 42480
rect 44730 42390 44760 42466
rect 44850 42210 44940 42480
rect 45180 41880 45300 42705
rect 46380 42690 46500 42810
rect 48060 42795 48180 42810
rect 46410 42480 46500 42690
rect 48060 42705 54434 42795
rect 48060 42690 48180 42705
rect 48090 42480 48180 42690
rect 45660 42466 45930 42480
rect 44610 41280 44730 41294
rect 44850 41866 44970 41880
rect 44850 41190 44970 41294
rect 45180 41280 45300 41310
rect 45420 41190 45540 41310
rect 45780 42390 45930 42466
rect 46320 42466 46560 42480
rect 45660 41280 45780 41294
rect 45900 42210 46050 42270
rect 45900 41340 45914 42210
rect 46036 41340 46050 42210
rect 45900 41280 46050 41340
rect 46320 41294 46380 42466
rect 46500 41294 46560 42466
rect 46980 42466 47220 42480
rect 46980 42390 47100 42466
rect 46320 41280 46560 41294
rect 46830 42210 46980 42270
rect 46830 41340 46844 42210
rect 46966 41340 46980 42210
rect 45930 41190 46050 41280
rect 46830 41190 46980 41340
rect 47100 41280 47220 41294
rect 47340 42466 47610 42480
rect 47460 42390 47610 42466
rect 48000 42466 48240 42480
rect 47340 41280 47460 41294
rect 47580 42210 47730 42270
rect 47580 41340 47594 42210
rect 47716 41340 47730 42210
rect 47580 41280 47730 41340
rect 48000 41294 48060 42466
rect 48180 41294 48240 42466
rect 48660 42466 48900 42480
rect 48660 42390 48780 42466
rect 48000 41280 48240 41294
rect 48510 42210 48660 42270
rect 48510 41340 48524 42210
rect 48646 41340 48660 42210
rect 47610 41190 47730 41280
rect 48510 41190 48660 41340
rect 48780 41280 48900 41294
rect 1155 41160 54240 41190
rect 1155 41040 1214 41160
rect 2086 41040 5220 41160
rect 5340 41040 5460 41160
rect 5580 41040 5700 41160
rect 5820 41040 5940 41160
rect 6060 41040 6180 41160
rect 6300 41040 6420 41160
rect 6540 41040 6660 41160
rect 6780 41040 6900 41160
rect 7020 41040 7140 41160
rect 7260 41040 7380 41160
rect 7500 41040 7620 41160
rect 7740 41040 7860 41160
rect 7980 41040 8100 41160
rect 8220 41040 8340 41160
rect 8460 41040 8580 41160
rect 8700 41040 8820 41160
rect 8940 41040 9060 41160
rect 9180 41040 9300 41160
rect 9420 41040 9540 41160
rect 9660 41040 9780 41160
rect 9900 41040 10020 41160
rect 10140 41040 10260 41160
rect 10380 41040 10500 41160
rect 10620 41040 10740 41160
rect 10860 41040 10980 41160
rect 11100 41040 11460 41160
rect 11580 41040 11700 41160
rect 11820 41040 11940 41160
rect 12060 41040 12180 41160
rect 12300 41040 12420 41160
rect 12540 41040 12900 41160
rect 13020 41040 13140 41160
rect 13260 41040 13380 41160
rect 13500 41040 13620 41160
rect 13740 41040 13860 41160
rect 13980 41040 14100 41160
rect 14220 41040 14340 41160
rect 14460 41040 14580 41160
rect 14700 41040 14820 41160
rect 14940 41040 15060 41160
rect 15180 41040 15300 41160
rect 15420 41040 15540 41160
rect 15660 41040 15780 41160
rect 15900 41040 16020 41160
rect 16140 41040 16260 41160
rect 16380 41040 16500 41160
rect 16620 41040 16740 41160
rect 16860 41040 16980 41160
rect 17100 41040 17220 41160
rect 17340 41040 17460 41160
rect 17580 41040 17940 41160
rect 18060 41040 18180 41160
rect 18300 41040 18420 41160
rect 18540 41040 18660 41160
rect 18780 41040 18900 41160
rect 19020 41040 19140 41160
rect 19260 41040 19380 41160
rect 19500 41040 19620 41160
rect 19740 41040 19860 41160
rect 19980 41040 20100 41160
rect 20220 41040 20340 41160
rect 20460 41040 20580 41160
rect 20700 41040 20820 41160
rect 20940 41040 21060 41160
rect 21180 41040 21540 41160
rect 21660 41040 21780 41160
rect 21900 41040 22020 41160
rect 22140 41040 22260 41160
rect 22380 41040 22500 41160
rect 22620 41040 22740 41160
rect 22860 41040 22980 41160
rect 23100 41040 23220 41160
rect 23340 41040 23460 41160
rect 23580 41040 23700 41160
rect 23820 41040 23940 41160
rect 24060 41040 24180 41160
rect 24300 41040 24420 41160
rect 24540 41040 24660 41160
rect 24780 41040 24900 41160
rect 25020 41040 25140 41160
rect 25260 41040 25380 41160
rect 25500 41040 25620 41160
rect 25740 41040 25860 41160
rect 25980 41040 26100 41160
rect 26220 41040 26340 41160
rect 26460 41040 26580 41160
rect 26700 41040 27060 41160
rect 27180 41040 27300 41160
rect 27420 41040 27540 41160
rect 27660 41040 27780 41160
rect 27900 41040 28260 41160
rect 28380 41040 28500 41160
rect 28620 41040 28740 41160
rect 28860 41040 28980 41160
rect 29100 41040 29220 41160
rect 29340 41040 29460 41160
rect 29580 41040 29700 41160
rect 29820 41040 29940 41160
rect 30060 41040 30180 41160
rect 30300 41040 30420 41160
rect 30540 41040 30660 41160
rect 30780 41040 31140 41160
rect 31260 41040 31380 41160
rect 31500 41040 31620 41160
rect 31740 41040 31860 41160
rect 31980 41040 32100 41160
rect 32220 41040 32580 41160
rect 32700 41040 32820 41160
rect 32940 41040 33060 41160
rect 33180 41040 33300 41160
rect 33420 41040 33780 41160
rect 33900 41040 34020 41160
rect 34140 41040 34260 41160
rect 34380 41040 34500 41160
rect 34620 41040 34740 41160
rect 34860 41040 34980 41160
rect 35100 41040 35220 41160
rect 35340 41040 35460 41160
rect 35580 41040 35700 41160
rect 35820 41040 35940 41160
rect 36060 41040 36180 41160
rect 36300 41040 36420 41160
rect 36540 41040 36660 41160
rect 36780 41040 36900 41160
rect 37020 41040 37140 41160
rect 37260 41040 37380 41160
rect 37500 41040 37620 41160
rect 37740 41040 37860 41160
rect 37980 41040 38100 41160
rect 38220 41040 38340 41160
rect 38460 41040 38580 41160
rect 38700 41040 38820 41160
rect 38940 41040 39060 41160
rect 39180 41040 39300 41160
rect 39420 41040 39540 41160
rect 39660 41040 39780 41160
rect 39900 41040 40020 41160
rect 40140 41040 40260 41160
rect 40380 41040 40500 41160
rect 40620 41040 40740 41160
rect 40860 41040 40980 41160
rect 41100 41040 41220 41160
rect 41340 41040 41460 41160
rect 41580 41040 41700 41160
rect 41820 41040 42180 41160
rect 42300 41040 42420 41160
rect 42540 41040 42660 41160
rect 42780 41040 42900 41160
rect 43020 41040 43380 41160
rect 43500 41040 43860 41160
rect 43980 41040 44100 41160
rect 44220 41040 44340 41160
rect 44460 41040 44580 41160
rect 44700 41040 45060 41160
rect 45180 41040 45300 41160
rect 45420 41040 45540 41160
rect 45660 41040 45780 41160
rect 45900 41040 46020 41160
rect 46140 41040 46260 41160
rect 46380 41040 46500 41160
rect 46620 41040 46740 41160
rect 46860 41040 46980 41160
rect 47100 41040 47220 41160
rect 47340 41040 47460 41160
rect 47580 41040 47700 41160
rect 47820 41040 47940 41160
rect 48060 41040 48180 41160
rect 48300 41040 48420 41160
rect 48540 41040 48660 41160
rect 48780 41040 48900 41160
rect 49020 41040 49140 41160
rect 49260 41040 49380 41160
rect 49500 41040 49620 41160
rect 49740 41040 49860 41160
rect 49980 41040 50100 41160
rect 50220 41040 53310 41160
rect 54180 41040 54240 41160
rect 1155 41010 54240 41040
rect 6060 40920 6180 41010
rect 5820 40876 5940 40920
rect 6300 40906 6420 40920
rect 5820 39810 5940 39854
rect 5820 39734 6300 39810
rect 5820 39720 6420 39734
rect 6540 40906 6660 40920
rect 8220 40906 8340 41010
rect 6660 40605 7260 40695
rect 8220 40320 8340 40334
rect 8460 40906 8580 40920
rect 8220 39795 8340 39810
rect 6540 39720 6660 39734
rect 5820 39495 5940 39510
rect 5700 39450 5940 39495
rect 6540 39510 6630 39720
rect 7035 39705 8340 39795
rect 5700 39420 6060 39450
rect 6300 39495 6660 39510
rect 7035 39495 7125 39705
rect 8220 39690 8340 39705
rect 6300 39420 7125 39495
rect 5700 39405 5940 39420
rect 5820 39390 5940 39405
rect 6060 39090 6180 39210
rect 6300 38880 6390 39420
rect 6540 39405 7125 39420
rect 6540 39390 6660 39405
rect 6540 38895 6660 38910
rect 6540 38805 7020 38895
rect 6540 38790 6660 38805
rect 8460 38880 8580 40334
rect 8700 40906 8820 41010
rect 8700 40320 8820 40334
rect 9660 40906 9780 41010
rect 9660 40320 9780 40334
rect 9900 40906 10020 40920
rect 9900 39495 10020 40334
rect 10140 40906 10260 41010
rect 11100 40920 11220 41010
rect 11850 40920 11970 41010
rect 10140 40320 10260 40334
rect 10620 40906 10740 40920
rect 10620 39720 10740 39734
rect 10860 40906 10980 40920
rect 11340 40876 11460 40920
rect 11340 39810 11460 39854
rect 10980 39734 11460 39810
rect 10860 39720 11460 39734
rect 11580 40906 11700 40920
rect 11820 40860 11970 40920
rect 11820 39990 11834 40860
rect 11956 39990 11970 40860
rect 11820 39930 11970 39990
rect 12240 40906 12480 40920
rect 11700 39734 11790 39810
rect 11580 39720 11790 39734
rect 12240 39734 12300 40906
rect 12420 39810 12480 40906
rect 12750 40860 12900 41010
rect 12750 39990 12764 40860
rect 12886 39990 12900 40860
rect 12750 39930 12900 39990
rect 13020 40906 13140 40920
rect 12420 39734 12540 39810
rect 12240 39720 12540 39734
rect 12900 39734 13020 39810
rect 13500 40906 13620 41010
rect 13500 40320 13620 40334
rect 13740 40906 13860 40920
rect 12900 39720 13140 39734
rect 10650 39510 10740 39720
rect 11820 39630 11910 39720
rect 9435 39405 10020 39495
rect 8700 39195 8820 39210
rect 9435 39195 9525 39405
rect 8700 39105 9525 39195
rect 8700 39090 8820 39105
rect 9900 38880 10020 39405
rect 10620 39420 10980 39510
rect 11820 39540 12210 39630
rect 12450 39510 12540 39720
rect 11220 39420 11340 39450
rect 10620 39390 10740 39420
rect 8430 38790 8580 38880
rect 5910 38190 6030 38280
rect 6540 38190 6660 38280
rect 8700 38190 8820 38280
rect 9900 38790 10050 38880
rect 10620 38895 10740 38910
rect 10500 38805 10740 38895
rect 10890 38880 10980 39420
rect 12450 39420 12660 39510
rect 12000 39330 12270 39420
rect 12180 39240 12270 39330
rect 12390 39390 12660 39420
rect 13020 39495 13140 39510
rect 13740 39495 13860 40334
rect 13980 40906 14100 41010
rect 13980 40320 14100 40334
rect 14460 40906 14580 40920
rect 14460 40320 14580 40334
rect 14700 40906 14820 41010
rect 14700 40320 14820 40334
rect 14940 40906 15060 40920
rect 14940 40320 15060 40334
rect 15180 40906 15300 41010
rect 15180 40320 15300 40334
rect 15660 40890 15780 41010
rect 15900 40890 16020 40920
rect 14460 40110 14550 40320
rect 14940 40230 15030 40320
rect 14670 40140 15030 40230
rect 14460 39990 14580 40110
rect 13020 39405 13860 39495
rect 13020 39390 13140 39405
rect 12390 39330 12540 39390
rect 11100 39195 11220 39210
rect 11100 39105 11580 39195
rect 11100 39090 11220 39105
rect 11820 39090 12090 39180
rect 12000 39030 12090 39090
rect 11580 38880 11790 38970
rect 12000 38940 12060 39030
rect 10620 38790 10740 38805
rect 12390 38820 12480 39330
rect 13020 39195 13140 39210
rect 13260 39195 13380 39210
rect 13020 39105 13380 39195
rect 13020 39090 13140 39105
rect 13260 39090 13380 39105
rect 12600 39030 12690 39090
rect 12900 38880 13140 38970
rect 13740 38880 13860 39405
rect 11820 38760 11970 38790
rect 11820 38280 11970 38310
rect 12240 38760 12480 38820
rect 12240 38340 12300 38760
rect 12420 38340 12480 38760
rect 12240 38280 12480 38340
rect 12750 38760 12900 38790
rect 9660 38190 9780 38280
rect 10620 38190 10740 38280
rect 11250 38190 11370 38280
rect 11850 38190 11970 38280
rect 12750 38190 12900 38310
rect 13740 38790 13890 38880
rect 14460 38670 14550 39990
rect 14670 39090 14760 40140
rect 14850 39795 15060 39810
rect 14850 39705 15660 39795
rect 14850 39690 15060 39705
rect 15900 39495 16020 40320
rect 16380 40906 16500 41010
rect 16380 39720 16500 39734
rect 16770 40906 16890 40920
rect 17010 40906 17130 41010
rect 17010 40320 17130 40334
rect 17670 40906 17790 41010
rect 17670 40320 17790 40334
rect 17910 40906 18030 40920
rect 17010 39810 17100 39990
rect 16890 39734 16920 39810
rect 16770 39720 16920 39734
rect 17010 39795 17220 39810
rect 17010 39720 17340 39795
rect 16620 39495 16740 39510
rect 15900 39405 16740 39495
rect 14760 39000 15090 39090
rect 15000 38970 15090 39000
rect 15000 38880 15270 38970
rect 14460 38580 14670 38670
rect 15660 38895 15780 38910
rect 15540 38805 15780 38895
rect 15660 38790 15780 38805
rect 15660 38550 15780 38580
rect 15900 38550 16020 39405
rect 16620 39390 16740 39405
rect 16830 39210 16920 39720
rect 17100 39705 17340 39720
rect 17100 39690 17220 39705
rect 17700 39720 17790 39990
rect 17880 39734 17910 39810
rect 17880 39720 18030 39734
rect 18300 40906 18420 41010
rect 18300 39720 18420 39734
rect 18540 40890 18660 40920
rect 18780 40890 18900 41010
rect 19260 40906 19380 41010
rect 17880 39210 17970 39720
rect 18060 39495 18180 39510
rect 18540 39495 18660 40320
rect 19260 39720 19380 39734
rect 19650 40906 19770 40920
rect 19890 40906 20010 41010
rect 19890 40320 20010 40334
rect 20940 40906 21060 41010
rect 20940 40320 21060 40334
rect 21180 40906 21300 40920
rect 19890 39810 19980 39990
rect 19770 39734 19800 39810
rect 19650 39720 19800 39734
rect 19890 39795 20100 39810
rect 19890 39720 20805 39795
rect 18060 39405 18660 39495
rect 18060 39390 18180 39405
rect 16380 39195 16500 39210
rect 16260 39180 16500 39195
rect 16260 39150 16620 39180
rect 16260 39105 16500 39150
rect 16380 39090 16500 39105
rect 16830 39090 17220 39210
rect 17580 39090 17970 39210
rect 18300 39180 18420 39210
rect 18180 39150 18420 39180
rect 16410 38880 16950 38940
rect 17100 38880 17190 39090
rect 17610 38880 17700 39090
rect 18300 39090 18420 39150
rect 17850 38880 18390 38940
rect 16500 38850 16860 38880
rect 16620 38730 16740 38760
rect 13500 38190 13620 38280
rect 14790 38190 14910 38280
rect 15660 38190 15780 38280
rect 16620 38190 16740 38310
rect 17940 38850 18300 38880
rect 18060 38730 18180 38760
rect 18060 38190 18180 38310
rect 18540 38550 18660 39405
rect 19500 39495 19620 39510
rect 18900 39405 19620 39495
rect 19500 39390 19620 39405
rect 19710 39210 19800 39720
rect 19980 39705 20805 39720
rect 19980 39690 20100 39705
rect 20715 39495 20805 39705
rect 21180 39495 21300 40334
rect 21420 40906 21540 41010
rect 22170 40920 22290 41010
rect 21420 40320 21540 40334
rect 21900 40906 22020 40920
rect 22140 40860 22290 40920
rect 22140 39990 22154 40860
rect 22276 39990 22290 40860
rect 22140 39930 22290 39990
rect 22560 40906 22800 40920
rect 22020 39734 22170 39810
rect 21900 39720 22170 39734
rect 22560 39734 22620 40906
rect 22740 39734 22800 40906
rect 23070 40860 23220 41010
rect 23070 39990 23084 40860
rect 23206 39990 23220 40860
rect 23070 39930 23220 39990
rect 23340 40906 23460 40920
rect 22560 39720 22800 39734
rect 23220 39734 23340 39810
rect 23220 39720 23460 39734
rect 23820 40890 23940 41010
rect 24210 40890 24330 40920
rect 24060 39720 24210 39840
rect 24780 40906 24900 41010
rect 24780 39720 24900 39734
rect 25170 40906 25290 40920
rect 25410 40906 25530 41010
rect 26460 40920 26580 41010
rect 25410 40320 25530 40334
rect 26220 40876 26340 40920
rect 25410 39810 25500 39990
rect 26700 40906 27300 40920
rect 26220 39810 26340 39854
rect 25290 39734 25320 39810
rect 25170 39720 25320 39734
rect 25410 39795 25620 39810
rect 25410 39720 25740 39795
rect 20715 39405 21300 39495
rect 18780 39195 18900 39210
rect 19260 39195 19380 39210
rect 18780 39180 19380 39195
rect 18780 39150 19500 39180
rect 18780 39105 19380 39150
rect 18780 39090 18900 39105
rect 19260 39090 19380 39105
rect 19710 39090 19740 39210
rect 19860 39090 20100 39210
rect 18780 38895 18900 38910
rect 18780 38805 19020 38895
rect 18780 38790 18900 38805
rect 19290 38880 19830 38940
rect 19980 38880 20070 39090
rect 21180 38880 21300 39405
rect 22650 39510 22740 39720
rect 22620 39390 22740 39510
rect 21540 39105 21660 39195
rect 22140 39150 22440 39240
rect 22650 39210 22740 39390
rect 24090 39210 24180 39720
rect 25020 39495 25140 39510
rect 24420 39405 25140 39495
rect 25020 39390 25140 39405
rect 25230 39210 25320 39720
rect 25500 39705 25740 39720
rect 25500 39690 25620 39705
rect 26220 39734 26700 39810
rect 26820 40830 27180 40906
rect 26220 39720 26820 39734
rect 27180 39720 27300 39734
rect 27900 40890 28020 40920
rect 28140 40890 28260 41010
rect 30540 40906 30660 41010
rect 30540 40320 30660 40334
rect 30780 40906 30900 40920
rect 26940 39630 27030 39720
rect 26730 39540 27030 39630
rect 26730 39510 26820 39540
rect 26340 39420 26460 39450
rect 26700 39390 26820 39510
rect 27180 39390 27300 39510
rect 22140 39120 22230 39150
rect 22650 39120 22800 39210
rect 21900 38880 22170 38970
rect 18780 38550 18900 38580
rect 19380 38850 19740 38880
rect 19500 38730 19620 38760
rect 18780 38190 18900 38280
rect 19500 38190 19620 38310
rect 21150 38790 21300 38880
rect 22710 38820 22800 39120
rect 23340 39195 23460 39210
rect 23820 39195 23940 39210
rect 23340 39105 23940 39195
rect 23340 39090 23460 39105
rect 23820 39090 23940 39105
rect 25230 39195 25620 39210
rect 26460 39195 26580 39210
rect 24900 39150 25020 39180
rect 22920 39030 23010 39090
rect 23220 38880 23460 38970
rect 22140 38760 22290 38790
rect 22140 38280 22290 38310
rect 22560 38760 22800 38820
rect 22560 38340 22620 38760
rect 22740 38340 22800 38760
rect 22560 38280 22800 38340
rect 23070 38760 23220 38790
rect 21420 38190 21540 38280
rect 22170 38190 22290 38280
rect 23070 38190 23220 38310
rect 23580 38895 23700 38910
rect 23820 38895 23940 38910
rect 23580 38805 23940 38895
rect 23580 38790 23700 38805
rect 23820 38790 23940 38805
rect 24090 38580 24180 39090
rect 25230 39105 26580 39195
rect 25230 39090 25620 39105
rect 26460 39090 26580 39105
rect 24810 38880 25350 38940
rect 25500 38880 25590 39090
rect 26730 38880 26820 39390
rect 26940 39210 27030 39270
rect 26940 39195 27060 39210
rect 27900 39195 28020 40320
rect 30540 39795 30660 39810
rect 29700 39705 30660 39795
rect 30540 39690 30660 39705
rect 30780 39795 30900 40334
rect 31020 40906 31140 41010
rect 31020 40320 31140 40334
rect 31980 40906 32100 41010
rect 31980 40320 32100 40334
rect 32220 40906 32340 40920
rect 31980 39795 32100 39810
rect 30780 39705 32100 39795
rect 26940 39105 28020 39195
rect 26940 39090 27060 39105
rect 24900 38850 25260 38880
rect 25020 38730 25140 38760
rect 23820 38190 23940 38280
rect 24300 38190 24420 38280
rect 25020 38190 25140 38310
rect 26670 38280 26730 38880
rect 26850 38280 26910 38880
rect 27900 38550 28020 39105
rect 28140 38790 28260 38910
rect 30780 38880 30900 39705
rect 31980 39690 32100 39705
rect 31020 39195 31140 39210
rect 31020 39105 31260 39195
rect 31020 39090 31140 39105
rect 32220 38880 32340 40334
rect 32460 40906 32580 41010
rect 33690 40920 33810 41010
rect 32460 40320 32580 40334
rect 33420 40906 33540 40920
rect 33660 40860 33810 40920
rect 33660 39990 33674 40860
rect 33796 39990 33810 40860
rect 33660 39930 33810 39990
rect 34080 40906 34320 40920
rect 33540 39734 33690 39810
rect 33420 39720 33690 39734
rect 34080 39734 34140 40906
rect 34260 39734 34320 40906
rect 34590 40860 34740 41010
rect 34590 39990 34604 40860
rect 34726 39990 34740 40860
rect 34590 39930 34740 39990
rect 34860 40906 34980 40920
rect 34080 39720 34320 39734
rect 34740 39734 34860 39810
rect 34740 39720 34980 39734
rect 36060 40906 36180 41010
rect 36060 39720 36180 39734
rect 36450 40906 36570 40920
rect 36690 40906 36810 41010
rect 36690 40320 36810 40334
rect 37740 40906 37860 41010
rect 37740 40320 37860 40334
rect 37980 40906 38100 40920
rect 36690 39810 36780 39990
rect 36570 39734 36600 39810
rect 36450 39720 36600 39734
rect 36690 39795 36900 39810
rect 36690 39720 37260 39795
rect 34170 39510 34260 39720
rect 34140 39390 34260 39510
rect 36300 39495 36420 39510
rect 35460 39405 36420 39495
rect 33420 39090 33540 39210
rect 33660 39150 33960 39240
rect 34170 39210 34260 39390
rect 33660 39120 33750 39150
rect 34170 39120 34320 39210
rect 33420 38880 33690 38970
rect 28140 38550 28260 38580
rect 30750 38790 30900 38880
rect 32190 38790 32340 38880
rect 34230 38820 34320 39120
rect 35595 39195 35685 39405
rect 36300 39390 36420 39405
rect 36510 39210 36600 39720
rect 36780 39705 37260 39720
rect 36780 39690 36900 39705
rect 37740 39795 37860 39810
rect 37380 39705 37860 39795
rect 37740 39690 37860 39705
rect 34980 39105 35685 39195
rect 36060 39180 36180 39210
rect 36060 39150 36300 39180
rect 36060 39090 36180 39150
rect 34440 39030 34530 39090
rect 36510 39090 36900 39210
rect 34740 38880 34980 38970
rect 36090 38880 36630 38940
rect 36780 38880 36870 39090
rect 37980 38880 38100 40334
rect 38220 40906 38340 41010
rect 38220 40320 38340 40334
rect 38940 40906 39060 41010
rect 38940 39720 39060 39734
rect 39330 40906 39450 40920
rect 39570 40906 39690 41010
rect 39570 40320 39690 40334
rect 40380 40906 40500 41010
rect 40380 40320 40500 40334
rect 40620 40906 40740 40920
rect 39570 39810 39660 39990
rect 39450 39734 39480 39810
rect 39330 39720 39480 39734
rect 39570 39795 39780 39810
rect 40620 39795 40740 40334
rect 40860 40906 40980 41010
rect 40860 40320 40980 40334
rect 41820 40890 41940 41010
rect 42060 40890 42180 40920
rect 39570 39720 40740 39795
rect 39180 39495 39300 39510
rect 38820 39405 39300 39495
rect 39180 39390 39300 39405
rect 39390 39210 39480 39720
rect 39660 39705 40740 39720
rect 39660 39690 39780 39705
rect 38940 39180 39060 39210
rect 38940 39150 39180 39180
rect 38940 39090 39060 39150
rect 39390 39090 39420 39210
rect 39540 39090 39780 39210
rect 39900 39195 40020 39210
rect 40380 39195 40500 39210
rect 39900 39105 40500 39195
rect 39900 39090 40020 39105
rect 40380 39090 40500 39105
rect 38970 38880 39510 38940
rect 39660 38880 39750 39090
rect 40620 38880 40740 39705
rect 42060 39495 42180 40320
rect 43020 40906 43140 41010
rect 43020 39720 43140 39734
rect 43410 40906 43530 40920
rect 43650 40906 43770 41010
rect 43650 40320 43770 40334
rect 44700 40890 44820 41010
rect 44940 40890 45060 40920
rect 45990 40906 46110 41010
rect 45990 40320 46110 40334
rect 46230 40906 46350 40920
rect 43530 39734 43560 39810
rect 43410 39720 43560 39734
rect 43650 39720 43740 39990
rect 43260 39495 43380 39510
rect 42060 39405 43380 39495
rect 33660 38760 33810 38790
rect 33660 38280 33810 38310
rect 34080 38760 34320 38820
rect 34080 38340 34140 38760
rect 34260 38340 34320 38760
rect 34080 38280 34320 38340
rect 34590 38760 34740 38790
rect 26280 38190 26400 38280
rect 27180 38190 27300 38280
rect 28140 38190 28260 38280
rect 31020 38190 31140 38280
rect 32460 38190 32580 38280
rect 33690 38190 33810 38280
rect 34590 38190 34740 38310
rect 36180 38850 36540 38880
rect 36300 38730 36420 38760
rect 36300 38190 36420 38310
rect 37500 38595 37620 38610
rect 36900 38505 37620 38595
rect 37500 38490 37620 38505
rect 37950 38790 38100 38880
rect 39060 38850 39420 38880
rect 39180 38730 39300 38760
rect 38220 38190 38340 38280
rect 39180 38190 39300 38310
rect 40620 38790 40770 38880
rect 41820 38895 41940 38910
rect 41700 38805 41940 38895
rect 41820 38790 41940 38805
rect 41820 38550 41940 38580
rect 42060 38550 42180 39405
rect 43260 39390 43380 39405
rect 43470 39210 43560 39720
rect 44940 39495 45060 40320
rect 46020 39810 46110 39990
rect 45900 39795 46110 39810
rect 45300 39720 46110 39795
rect 46200 39734 46230 39810
rect 46200 39720 46350 39734
rect 46620 40906 46740 41010
rect 46620 39720 46740 39734
rect 47580 40906 47700 41010
rect 47580 39720 47700 39734
rect 47970 40906 48090 40920
rect 48210 40906 48330 41010
rect 48210 40320 48330 40334
rect 49260 40906 49380 41010
rect 49260 40320 49380 40334
rect 49500 40906 49620 40920
rect 48210 39810 48300 39990
rect 48090 39734 48120 39810
rect 47970 39720 48120 39734
rect 48210 39795 48420 39810
rect 48210 39720 49125 39795
rect 45300 39705 46020 39720
rect 45900 39690 46020 39705
rect 45900 39495 46020 39510
rect 44940 39405 46020 39495
rect 43020 39195 43140 39210
rect 42660 39180 43140 39195
rect 43470 39195 43860 39210
rect 42660 39150 43260 39180
rect 42660 39105 43140 39150
rect 43020 39090 43140 39105
rect 43470 39105 43980 39195
rect 43470 39090 43860 39105
rect 43050 38880 43590 38940
rect 43740 38880 43830 39090
rect 43140 38850 43500 38880
rect 43260 38730 43380 38760
rect 40380 38190 40500 38280
rect 41820 38190 41940 38280
rect 43260 38190 43380 38310
rect 44700 38550 44820 38580
rect 44940 38550 45060 39405
rect 45900 39390 46020 39405
rect 46200 39210 46290 39720
rect 46380 39390 46500 39510
rect 46740 39405 47820 39495
rect 48030 39210 48120 39720
rect 48300 39705 49125 39720
rect 48300 39690 48420 39705
rect 49035 39495 49125 39705
rect 49260 39690 49380 39810
rect 49500 39495 49620 40334
rect 49740 40906 49860 41010
rect 49740 40320 49860 40334
rect 49035 39405 49620 39495
rect 45900 39090 46140 39210
rect 46260 39090 46290 39210
rect 46620 39195 46740 39210
rect 46620 39180 46860 39195
rect 46500 39150 46860 39180
rect 45930 38880 46020 39090
rect 46620 39105 46860 39150
rect 46620 39090 46740 39105
rect 47580 39195 47700 39210
rect 46980 39180 47700 39195
rect 46980 39150 47820 39180
rect 46980 39105 47700 39150
rect 47580 39090 47700 39105
rect 48030 39090 48420 39210
rect 46170 38880 46710 38940
rect 47610 38880 48150 38940
rect 48300 38880 48390 39090
rect 49500 38880 49620 39405
rect 45420 38595 45540 38610
rect 45420 38505 45900 38595
rect 45420 38490 45540 38505
rect 46260 38850 46620 38880
rect 46380 38730 46500 38760
rect 44700 38190 44820 38280
rect 46380 38190 46500 38310
rect 47700 38850 48060 38880
rect 47820 38730 47940 38760
rect 47820 38190 47940 38310
rect 49470 38790 49620 38880
rect 49740 38190 49860 38280
rect 3135 38160 52260 38190
rect 3135 38040 3194 38160
rect 4066 38040 5220 38160
rect 5340 38040 5460 38160
rect 5580 38040 5700 38160
rect 5820 38040 6180 38160
rect 6300 38040 6420 38160
rect 6540 38040 6660 38160
rect 6780 38040 6900 38160
rect 7020 38040 7140 38160
rect 7260 38040 7380 38160
rect 7500 38040 7620 38160
rect 7740 38040 7860 38160
rect 7980 38040 8100 38160
rect 8220 38040 8340 38160
rect 8460 38040 8580 38160
rect 8700 38040 8820 38160
rect 8940 38040 9060 38160
rect 9180 38040 9300 38160
rect 9420 38040 9540 38160
rect 9660 38040 9780 38160
rect 9900 38040 10020 38160
rect 10140 38040 10260 38160
rect 10380 38040 10500 38160
rect 10620 38040 10740 38160
rect 10860 38040 10980 38160
rect 11100 38040 11220 38160
rect 11340 38040 11460 38160
rect 11580 38040 11700 38160
rect 11820 38040 11940 38160
rect 12060 38040 12420 38160
rect 12540 38040 12900 38160
rect 13020 38040 13140 38160
rect 13260 38040 13380 38160
rect 13500 38040 13620 38160
rect 13740 38040 13860 38160
rect 13980 38040 14100 38160
rect 14220 38040 14340 38160
rect 14460 38040 14580 38160
rect 14700 38040 14820 38160
rect 14940 38040 15300 38160
rect 15420 38040 15540 38160
rect 15660 38040 15780 38160
rect 15900 38040 16020 38160
rect 16140 38040 16260 38160
rect 16380 38040 16500 38160
rect 16620 38040 16740 38160
rect 16860 38040 16980 38160
rect 17100 38040 17220 38160
rect 17340 38040 17460 38160
rect 17580 38040 17700 38160
rect 17820 38040 17940 38160
rect 18060 38040 18420 38160
rect 18540 38040 18660 38160
rect 18780 38040 18900 38160
rect 19020 38040 19140 38160
rect 19260 38040 19380 38160
rect 19500 38040 19620 38160
rect 19740 38040 19860 38160
rect 19980 38040 20100 38160
rect 20220 38040 20340 38160
rect 20460 38040 20580 38160
rect 20700 38040 20820 38160
rect 20940 38040 21060 38160
rect 21180 38040 21300 38160
rect 21420 38040 21540 38160
rect 21660 38040 21780 38160
rect 21900 38040 22020 38160
rect 22140 38040 22260 38160
rect 22380 38040 22740 38160
rect 22860 38040 22980 38160
rect 23100 38040 23220 38160
rect 23340 38040 23460 38160
rect 23580 38040 23700 38160
rect 23820 38040 24180 38160
rect 24300 38040 24420 38160
rect 24540 38040 24660 38160
rect 24780 38040 24900 38160
rect 25020 38040 25140 38160
rect 25260 38040 25620 38160
rect 25740 38040 25860 38160
rect 25980 38040 26100 38160
rect 26220 38040 26340 38160
rect 26460 38040 26580 38160
rect 26700 38040 26820 38160
rect 26940 38040 27060 38160
rect 27180 38040 27300 38160
rect 27420 38040 27540 38160
rect 27660 38040 27780 38160
rect 27900 38040 28260 38160
rect 28380 38040 28500 38160
rect 28620 38040 28740 38160
rect 28860 38040 28980 38160
rect 29100 38040 29220 38160
rect 29340 38040 29460 38160
rect 29580 38040 29700 38160
rect 29820 38040 29940 38160
rect 30060 38040 30180 38160
rect 30300 38040 30420 38160
rect 30540 38040 30660 38160
rect 30780 38040 30900 38160
rect 31020 38040 31140 38160
rect 31260 38040 31380 38160
rect 31500 38040 31620 38160
rect 31740 38040 31860 38160
rect 31980 38040 32100 38160
rect 32220 38040 32340 38160
rect 32460 38040 32580 38160
rect 32700 38040 32820 38160
rect 32940 38040 33060 38160
rect 33180 38040 33300 38160
rect 33420 38040 33780 38160
rect 33900 38040 34020 38160
rect 34140 38040 34260 38160
rect 34380 38040 34500 38160
rect 34620 38040 34740 38160
rect 34860 38040 34980 38160
rect 35100 38040 35220 38160
rect 35340 38040 35460 38160
rect 35580 38040 35700 38160
rect 35820 38040 35940 38160
rect 36060 38040 36180 38160
rect 36300 38040 36420 38160
rect 36540 38040 36660 38160
rect 36780 38040 36900 38160
rect 37020 38040 37140 38160
rect 37260 38040 37380 38160
rect 37500 38040 37620 38160
rect 37740 38040 37860 38160
rect 37980 38040 38100 38160
rect 38220 38040 38340 38160
rect 38460 38040 38580 38160
rect 38700 38040 38820 38160
rect 38940 38040 39300 38160
rect 39420 38040 39540 38160
rect 39660 38040 39780 38160
rect 39900 38040 40020 38160
rect 40140 38040 40260 38160
rect 40380 38040 40500 38160
rect 40620 38040 40740 38160
rect 40860 38040 40980 38160
rect 41100 38040 41220 38160
rect 41340 38040 41460 38160
rect 41580 38040 41700 38160
rect 41820 38040 41940 38160
rect 42060 38040 42180 38160
rect 42300 38040 42420 38160
rect 42540 38040 42660 38160
rect 42780 38040 42900 38160
rect 43020 38040 43140 38160
rect 43260 38040 43380 38160
rect 43500 38040 43860 38160
rect 43980 38040 44100 38160
rect 44220 38040 44340 38160
rect 44460 38040 44580 38160
rect 44700 38040 44820 38160
rect 44940 38040 45060 38160
rect 45180 38040 45300 38160
rect 45420 38040 45540 38160
rect 45660 38040 45780 38160
rect 45900 38040 46020 38160
rect 46140 38040 46260 38160
rect 46380 38040 46500 38160
rect 46620 38040 46740 38160
rect 46860 38040 46980 38160
rect 47100 38040 47220 38160
rect 47340 38040 47460 38160
rect 47580 38040 47940 38160
rect 48060 38040 48420 38160
rect 48540 38040 48660 38160
rect 48780 38040 48900 38160
rect 49020 38040 49140 38160
rect 49260 38040 49380 38160
rect 49500 38040 49860 38160
rect 49980 38040 50100 38160
rect 50220 38040 51330 38160
rect 52200 38040 52260 38160
rect 3135 38010 52260 38040
rect 6060 37920 6180 38010
rect 7260 37920 7380 38010
rect 5790 37320 5940 37410
rect 7020 37890 7140 37920
rect 7020 37710 7140 37740
rect 7260 37620 7380 37650
rect 7620 37605 8220 37695
rect 5580 36390 5700 36510
rect 5580 35866 5700 35880
rect 5580 35190 5700 35294
rect 5820 35866 5940 37320
rect 6060 37095 6180 37110
rect 6780 37095 6900 37110
rect 6060 37005 6900 37095
rect 6060 36990 6180 37005
rect 6780 36990 6900 37005
rect 7020 35880 7140 37590
rect 7260 37395 7380 37410
rect 7260 37305 7500 37395
rect 7260 37290 7380 37305
rect 8700 37890 8820 38010
rect 10860 37920 10980 38010
rect 8700 37440 8820 37470
rect 8580 37320 8940 37350
rect 11100 37320 11250 37410
rect 12540 37890 12660 38010
rect 12540 37440 12660 37470
rect 12420 37320 12780 37350
rect 13620 37605 14940 37695
rect 15420 37890 15540 38010
rect 16950 37920 17070 38010
rect 18060 37920 18180 38010
rect 19500 37920 19620 38010
rect 20940 37920 21060 38010
rect 22380 37920 22500 38010
rect 23820 37920 23940 38010
rect 25500 37920 25620 38010
rect 15420 37440 15540 37470
rect 15300 37320 15660 37350
rect 16620 37530 16830 37620
rect 8250 37110 8340 37320
rect 8490 37260 9030 37320
rect 8220 36990 8460 37110
rect 8580 36990 8610 37110
rect 8940 37095 9060 37110
rect 10860 37095 10980 37110
rect 8940 37050 10980 37095
rect 8820 37020 10980 37050
rect 8940 37005 10980 37020
rect 8940 36990 9060 37005
rect 10860 36990 10980 37005
rect 8220 36480 8340 36510
rect 8520 36480 8610 36990
rect 8700 36795 8820 36810
rect 10860 36795 10980 36810
rect 8700 36705 10980 36795
rect 8700 36690 8820 36705
rect 10860 36690 10980 36705
rect 9180 36495 9300 36510
rect 11100 36495 11220 37320
rect 12090 37110 12180 37320
rect 12330 37260 12870 37320
rect 12060 36990 12450 37110
rect 14970 37110 15060 37320
rect 15210 37260 15750 37320
rect 12780 37095 12900 37110
rect 14700 37095 14820 37110
rect 12780 37050 14820 37095
rect 12660 37020 14820 37050
rect 12780 37005 14820 37020
rect 12780 36990 12900 37005
rect 14700 36990 14820 37005
rect 14940 36990 15330 37110
rect 15660 37095 15780 37110
rect 15660 37050 15900 37095
rect 15540 37020 15900 37050
rect 15660 37005 15900 37020
rect 15660 36990 15780 37005
rect 8220 36390 8430 36480
rect 8520 36466 8670 36480
rect 8520 36390 8550 36466
rect 8340 36210 8430 36390
rect 5820 35280 5940 35294
rect 6060 35866 6180 35880
rect 6060 35190 6180 35294
rect 7020 35280 7140 35310
rect 7260 35190 7380 35310
rect 8310 35866 8430 35880
rect 8310 35190 8430 35294
rect 8550 35280 8670 35294
rect 8940 36466 9060 36480
rect 9180 36405 11220 36495
rect 9180 36390 9300 36405
rect 8940 35190 9060 35294
rect 10860 35866 10980 35880
rect 10860 35190 10980 35294
rect 11100 35866 11220 36405
rect 11460 36405 11820 36495
rect 12360 36480 12450 36990
rect 12540 36795 12660 36810
rect 12540 36705 13740 36795
rect 12540 36690 12660 36705
rect 12180 36210 12270 36480
rect 12360 36466 12510 36480
rect 12360 36390 12390 36466
rect 11100 35280 11220 35294
rect 11340 35866 11460 35880
rect 11340 35190 11460 35294
rect 12150 35866 12270 35880
rect 12150 35190 12270 35294
rect 12390 35280 12510 35294
rect 12780 36466 12900 36480
rect 14940 36495 15060 36510
rect 13140 36480 15060 36495
rect 15240 36480 15330 36990
rect 15420 36795 15540 36810
rect 15420 36705 15660 36795
rect 15420 36690 15540 36705
rect 13140 36405 15150 36480
rect 14940 36390 15150 36405
rect 15240 36466 15390 36480
rect 15240 36390 15270 36466
rect 15060 36210 15150 36390
rect 12780 35190 12900 35294
rect 15030 35866 15150 35880
rect 15030 35190 15150 35294
rect 15270 35280 15390 35294
rect 15660 36466 15780 36480
rect 16620 36210 16710 37530
rect 18300 37320 18450 37410
rect 19740 37320 19890 37410
rect 17160 37230 17430 37320
rect 17160 37200 17250 37230
rect 16920 37110 17250 37200
rect 16140 36195 16260 36210
rect 16620 36195 16740 36210
rect 16140 36105 16740 36195
rect 16140 36090 16260 36105
rect 16620 36090 16740 36105
rect 15660 35190 15780 35294
rect 16620 35880 16710 36090
rect 16830 36060 16920 37110
rect 18060 37095 18180 37110
rect 17700 37005 18180 37095
rect 18060 36990 18180 37005
rect 17010 36390 17100 36510
rect 17220 36405 17820 36495
rect 16830 35970 17190 36060
rect 17100 35880 17190 35970
rect 16620 35866 16740 35880
rect 16620 35280 16740 35294
rect 16860 35866 16980 35880
rect 16860 35190 16980 35294
rect 17100 35866 17220 35880
rect 17100 35280 17220 35294
rect 17340 35866 17460 35880
rect 17340 35190 17460 35294
rect 18060 35866 18180 35880
rect 18060 35190 18180 35294
rect 18300 35866 18420 37320
rect 19740 36495 19860 37320
rect 21300 37320 21330 37410
rect 22620 37320 22770 37410
rect 23820 37620 23940 37650
rect 22890 37320 23820 37395
rect 20940 36990 21060 37110
rect 18660 36405 19860 36495
rect 18300 35280 18420 35294
rect 18540 35866 18660 35880
rect 18540 35190 18660 35294
rect 19500 35866 19620 35880
rect 19500 35190 19620 35294
rect 19740 35866 19860 36405
rect 19980 36390 20100 36510
rect 19740 35280 19860 35294
rect 19980 35866 20100 35880
rect 19980 35190 20100 35294
rect 20940 35866 21060 35880
rect 20940 35190 21060 35294
rect 21180 35866 21300 37290
rect 22620 37305 23820 37320
rect 21420 37095 21540 37110
rect 21420 37005 22380 37095
rect 21420 36990 21540 37005
rect 21420 36390 21540 36510
rect 21180 35280 21300 35294
rect 21420 35866 21540 35880
rect 21420 35190 21540 35294
rect 22380 35866 22500 35880
rect 22380 35190 22500 35294
rect 22620 35866 22740 37305
rect 24060 35880 24180 37650
rect 25230 37320 25380 37410
rect 26700 37890 26820 38010
rect 27900 37920 28020 38010
rect 29100 37920 29220 38010
rect 26700 37440 26820 37470
rect 26580 37320 26940 37350
rect 28140 37320 28290 37410
rect 29340 37320 29490 37410
rect 30300 37890 30420 38010
rect 31260 37920 31380 38010
rect 30300 37440 30420 37470
rect 30180 37320 30540 37350
rect 31260 37620 31380 37650
rect 31020 37395 31140 37410
rect 31260 37395 31380 37410
rect 25260 36495 25380 37320
rect 26490 37260 27030 37320
rect 25740 37095 25860 37110
rect 26460 37095 26580 37110
rect 25740 37050 26580 37095
rect 27180 37110 27270 37320
rect 25740 37020 26700 37050
rect 26910 37095 27300 37110
rect 25740 37005 26580 37020
rect 25740 36990 25860 37005
rect 26460 36990 26580 37005
rect 26910 37005 27420 37095
rect 26910 36990 27300 37005
rect 27900 36990 28020 37110
rect 26700 36795 26820 36810
rect 25620 36705 26820 36795
rect 26700 36690 26820 36705
rect 26220 36495 26340 36510
rect 25260 36405 26340 36495
rect 26910 36480 27000 36990
rect 28140 36795 28260 37320
rect 28380 37095 28500 37110
rect 28380 37005 29100 37095
rect 28380 36990 28500 37005
rect 29340 37095 29460 37320
rect 30090 37260 30630 37320
rect 29340 37005 30060 37095
rect 27300 36705 28260 36795
rect 27180 36480 27300 36510
rect 22620 35280 22740 35294
rect 22860 35866 22980 35880
rect 22860 35190 22980 35294
rect 23820 35190 23940 35310
rect 24060 35280 24180 35310
rect 25020 35866 25140 35880
rect 25020 35190 25140 35294
rect 25260 35866 25380 36405
rect 26220 36390 26340 36405
rect 26460 36466 26580 36480
rect 25260 35280 25380 35294
rect 25500 35866 25620 35880
rect 25500 35190 25620 35294
rect 26460 35190 26580 35294
rect 26850 36466 27000 36480
rect 26970 36390 27000 36466
rect 27090 36390 27300 36480
rect 27090 36210 27180 36390
rect 26850 35280 26970 35294
rect 27090 35866 27210 35880
rect 27090 35190 27210 35294
rect 27900 35866 28020 35880
rect 27900 35190 28020 35294
rect 28140 35866 28260 36705
rect 28380 36495 28500 36510
rect 28380 36405 28860 36495
rect 28380 36390 28500 36405
rect 28140 35280 28260 35294
rect 28380 35866 28500 35880
rect 28380 35190 28500 35294
rect 29100 35866 29220 35880
rect 29100 35190 29220 35294
rect 29340 35866 29460 37005
rect 30780 37110 30870 37320
rect 31020 37305 31380 37395
rect 31020 37290 31140 37305
rect 31260 37290 31380 37305
rect 30180 37020 30300 37050
rect 30510 36990 30900 37110
rect 30510 36480 30600 36990
rect 31500 36795 31620 37650
rect 32460 37890 32580 38010
rect 33660 37920 33780 38010
rect 32460 37440 32580 37470
rect 32340 37320 32700 37350
rect 32010 37110 32100 37320
rect 32250 37260 32790 37320
rect 33060 37320 33270 37395
rect 33390 37320 33540 37410
rect 34620 37920 34740 38010
rect 33060 37305 33540 37320
rect 31980 37095 32370 37110
rect 31860 37005 32370 37095
rect 32580 37020 32700 37050
rect 31980 36990 32370 37005
rect 31980 36795 32100 36810
rect 31500 36705 32100 36795
rect 30780 36495 30900 36510
rect 31260 36495 31380 36510
rect 30780 36480 31380 36495
rect 30060 36466 30180 36480
rect 29340 35280 29460 35294
rect 29580 35866 29700 35880
rect 29580 35190 29700 35294
rect 30060 35190 30180 35294
rect 30450 36466 30600 36480
rect 30570 36390 30600 36466
rect 30690 36405 31380 36480
rect 30690 36390 30900 36405
rect 31260 36390 31380 36405
rect 30690 36210 30780 36390
rect 31500 35880 31620 36705
rect 31980 36690 32100 36705
rect 32280 36480 32370 36990
rect 32460 36690 32580 36810
rect 32100 36210 32190 36480
rect 32280 36466 32430 36480
rect 32280 36390 32310 36466
rect 30450 35280 30570 35294
rect 30690 35866 30810 35880
rect 30690 35190 30810 35294
rect 31260 35190 31380 35310
rect 31500 35280 31620 35310
rect 32070 35866 32190 35880
rect 32070 35190 32190 35294
rect 32310 35280 32430 35294
rect 32700 36466 32820 36480
rect 33180 36390 33300 36510
rect 32700 35190 32820 35294
rect 33180 35866 33300 35880
rect 33180 35190 33300 35294
rect 33420 35866 33540 37305
rect 34980 37320 35010 37410
rect 35820 37890 35970 38010
rect 36750 37920 36870 38010
rect 38940 37920 39060 38010
rect 39900 37920 40020 38010
rect 35820 37410 35970 37440
rect 36240 37860 36480 37920
rect 36240 37440 36300 37860
rect 36420 37440 36480 37860
rect 36240 37380 36480 37440
rect 36750 37890 36900 37920
rect 36750 37410 36900 37440
rect 33660 37095 33780 37110
rect 33660 37005 34380 37095
rect 33660 36990 33780 37005
rect 33420 35280 33540 35294
rect 33660 35866 33780 35880
rect 33660 35190 33780 35294
rect 34620 35866 34740 35880
rect 34620 35190 34740 35294
rect 34860 35866 34980 37290
rect 35580 37230 35820 37320
rect 36030 37110 36120 37170
rect 35100 37095 35220 37110
rect 35580 37095 35700 37110
rect 35100 37005 35700 37095
rect 35100 36990 35220 37005
rect 35580 36990 35700 37005
rect 36240 37080 36330 37380
rect 38940 37620 39060 37650
rect 36870 37230 37140 37320
rect 38940 37395 39060 37410
rect 37380 37305 39060 37395
rect 38940 37290 39060 37305
rect 36240 36990 36390 37080
rect 36810 37050 36900 37080
rect 36300 36810 36390 36990
rect 36600 36960 36900 37050
rect 39180 37095 39300 37650
rect 40290 37868 40530 37920
rect 40290 37746 40350 37868
rect 40470 37746 40530 37868
rect 40290 37710 40530 37746
rect 40290 37590 40350 37710
rect 40470 37590 40530 37710
rect 40290 37522 40530 37590
rect 40290 37402 40350 37522
rect 40470 37402 40530 37522
rect 40290 37320 40530 37402
rect 40800 37906 40920 38010
rect 41580 37920 41700 38010
rect 41580 37620 41700 37650
rect 40800 37320 40920 37334
rect 40140 37095 40260 37110
rect 39180 37005 40260 37095
rect 36300 36690 36420 36810
rect 36300 36480 36390 36690
rect 35580 36466 35820 36480
rect 34860 35280 34980 35294
rect 35100 35866 35220 35880
rect 35100 35190 35220 35294
rect 35700 36390 35820 36466
rect 36240 36466 36480 36480
rect 35580 35280 35700 35294
rect 35820 36210 35970 36270
rect 35820 35340 35834 36210
rect 35956 35340 35970 36210
rect 35820 35190 35970 35340
rect 36240 35294 36300 36466
rect 36420 35294 36480 36466
rect 36870 36466 37140 36480
rect 36870 36390 37020 36466
rect 36240 35280 36480 35294
rect 36750 36210 36900 36270
rect 36750 35340 36764 36210
rect 36886 35340 36900 36210
rect 36750 35280 36900 35340
rect 39180 35880 39300 37005
rect 40140 36990 40260 37005
rect 40170 36930 40260 36990
rect 40380 36810 40470 37320
rect 41580 37395 41700 37410
rect 41220 37305 41700 37395
rect 41580 37290 41700 37305
rect 39900 36795 40020 36810
rect 39540 36705 40020 36795
rect 39900 36690 40020 36705
rect 40380 36690 40500 36810
rect 40740 36750 40860 36780
rect 40380 36660 40470 36690
rect 40170 36570 40470 36660
rect 41820 36795 41940 37650
rect 42300 37906 42420 37920
rect 42300 37320 42420 37334
rect 42540 37906 42660 37920
rect 42780 37890 42900 38010
rect 43740 37920 43860 38010
rect 42780 37440 42900 37470
rect 43020 37906 43140 37920
rect 42660 37334 43020 37350
rect 42540 37320 43140 37334
rect 42330 37110 42420 37320
rect 42570 37260 43110 37320
rect 42300 37095 42690 37110
rect 42180 37005 42690 37095
rect 43020 37095 43140 37110
rect 43260 37095 43380 37110
rect 43020 37050 43380 37095
rect 42900 37020 43380 37050
rect 42300 36990 42690 37005
rect 43020 37005 43380 37020
rect 43020 36990 43140 37005
rect 43260 36990 43380 37005
rect 42300 36795 42420 36810
rect 41820 36705 42420 36795
rect 40170 36480 40260 36570
rect 37020 35280 37140 35294
rect 36750 35190 36870 35280
rect 38940 35190 39060 35310
rect 39180 35280 39300 35310
rect 39900 36466 40020 36480
rect 40380 36466 40980 36480
rect 40020 35294 40380 35370
rect 40500 36390 40980 36466
rect 40860 36346 40980 36390
rect 39900 35280 40500 35294
rect 41820 35880 41940 36705
rect 42300 36690 42420 36705
rect 42600 36480 42690 36990
rect 42780 36690 42900 36810
rect 42420 36210 42510 36480
rect 42600 36466 42750 36480
rect 42600 36390 42630 36466
rect 40860 35280 40980 35324
rect 40620 35190 40740 35280
rect 41580 35190 41700 35310
rect 41820 35280 41940 35310
rect 42390 35866 42510 35880
rect 42390 35190 42510 35294
rect 42630 35280 42750 35294
rect 43020 36466 43140 36480
rect 43500 35880 43620 37650
rect 43740 37620 43860 37650
rect 44460 37906 44580 37920
rect 44700 37890 44820 38010
rect 44700 37440 44820 37470
rect 44940 37906 45060 37920
rect 44580 37334 44940 37350
rect 44460 37320 45060 37334
rect 45180 37906 45300 37920
rect 45180 37320 45300 37334
rect 46140 37906 46260 38010
rect 46530 37906 46650 37920
rect 46140 37320 46260 37334
rect 46380 37334 46530 37410
rect 46380 37320 46650 37334
rect 47580 37906 47700 37920
rect 47820 37890 47940 38010
rect 47820 37440 47940 37470
rect 48060 37906 48180 37920
rect 47700 37334 48060 37350
rect 47580 37320 48180 37334
rect 48300 37906 48420 37920
rect 48300 37320 48420 37334
rect 49350 37906 49470 37920
rect 49740 37906 49860 38010
rect 49470 37334 49620 37410
rect 49350 37320 49620 37334
rect 49740 37320 49860 37334
rect 44490 37260 45030 37320
rect 44460 37095 44580 37110
rect 44100 37050 44580 37095
rect 45180 37110 45270 37320
rect 44100 37020 44700 37050
rect 44100 37005 44580 37020
rect 44460 36990 44580 37005
rect 44910 36990 45300 37110
rect 45420 37095 45540 37110
rect 46140 37095 46260 37110
rect 45420 37005 46260 37095
rect 45420 36990 45540 37005
rect 46140 36990 46260 37005
rect 44910 36480 45000 36990
rect 45180 36495 45300 36510
rect 46380 36495 46500 37320
rect 47610 37260 48150 37320
rect 48300 37110 48390 37320
rect 47700 37020 47820 37050
rect 48030 36990 48420 37110
rect 47820 36690 47940 36810
rect 45180 36480 46500 36495
rect 44460 36466 44580 36480
rect 43260 35595 43380 35610
rect 43260 35505 43500 35595
rect 43260 35490 43380 35505
rect 43020 35190 43140 35294
rect 43500 35280 43620 35310
rect 43740 35190 43860 35310
rect 44460 35190 44580 35294
rect 44850 36466 45000 36480
rect 44970 36390 45000 36466
rect 45090 36405 46500 36480
rect 45090 36390 45300 36405
rect 45090 36210 45180 36390
rect 44850 35280 44970 35294
rect 45090 35866 45210 35880
rect 45090 35190 45210 35294
rect 46140 35866 46260 35880
rect 46140 35190 46260 35294
rect 46380 35866 46500 36405
rect 48030 36480 48120 36990
rect 49500 36795 49620 37320
rect 49035 36705 49620 36795
rect 48300 36495 48420 36510
rect 49035 36495 49125 36705
rect 48300 36480 49125 36495
rect 47580 36466 47700 36480
rect 46380 35280 46500 35294
rect 46620 35866 46740 35880
rect 46620 35190 46740 35294
rect 47580 35190 47700 35294
rect 47970 36466 48120 36480
rect 48090 36390 48120 36466
rect 48210 36405 49125 36480
rect 48210 36390 48420 36405
rect 49260 36390 49380 36510
rect 48210 36210 48300 36390
rect 47970 35280 48090 35294
rect 48210 35866 48330 35880
rect 48210 35190 48330 35294
rect 49260 35866 49380 35880
rect 49260 35190 49380 35294
rect 49500 35866 49620 36705
rect 49500 35280 49620 35294
rect 49740 35866 49860 35880
rect 49740 35190 49860 35294
rect 1155 35160 54240 35190
rect 1155 35040 1214 35160
rect 2086 35040 5220 35160
rect 5340 35040 5460 35160
rect 5580 35040 5700 35160
rect 5820 35040 5940 35160
rect 6060 35040 6180 35160
rect 6300 35040 6420 35160
rect 6540 35040 6660 35160
rect 6780 35040 6900 35160
rect 7020 35040 7380 35160
rect 7500 35040 7620 35160
rect 7740 35040 7860 35160
rect 7980 35040 8100 35160
rect 8220 35040 8580 35160
rect 8700 35040 8820 35160
rect 8940 35040 9060 35160
rect 9180 35040 9300 35160
rect 9420 35040 9540 35160
rect 9660 35040 9780 35160
rect 9900 35040 10020 35160
rect 10140 35040 10260 35160
rect 10380 35040 10500 35160
rect 10620 35040 10740 35160
rect 10860 35040 10980 35160
rect 11100 35040 11220 35160
rect 11340 35040 11460 35160
rect 11580 35040 11700 35160
rect 11820 35040 11940 35160
rect 12060 35040 12420 35160
rect 12540 35040 12660 35160
rect 12780 35040 12900 35160
rect 13020 35040 13140 35160
rect 13260 35040 13380 35160
rect 13500 35040 13620 35160
rect 13740 35040 13860 35160
rect 13980 35040 14100 35160
rect 14220 35040 14340 35160
rect 14460 35040 14580 35160
rect 14700 35040 14820 35160
rect 14940 35040 15060 35160
rect 15180 35040 15300 35160
rect 15420 35040 15540 35160
rect 15660 35040 15780 35160
rect 15900 35040 16020 35160
rect 16140 35040 16260 35160
rect 16380 35040 16500 35160
rect 16620 35040 16980 35160
rect 17100 35040 17460 35160
rect 17580 35040 17700 35160
rect 17820 35040 17940 35160
rect 18060 35040 18180 35160
rect 18300 35040 18420 35160
rect 18540 35040 18660 35160
rect 18780 35040 18900 35160
rect 19020 35040 19140 35160
rect 19260 35040 19380 35160
rect 19500 35040 19860 35160
rect 19980 35040 20100 35160
rect 20220 35040 20340 35160
rect 20460 35040 20580 35160
rect 20700 35040 20820 35160
rect 20940 35040 21060 35160
rect 21180 35040 21300 35160
rect 21420 35040 21540 35160
rect 21660 35040 21780 35160
rect 21900 35040 22020 35160
rect 22140 35040 22260 35160
rect 22380 35040 22500 35160
rect 22620 35040 22740 35160
rect 22860 35040 22980 35160
rect 23100 35040 23220 35160
rect 23340 35040 23460 35160
rect 23580 35040 23700 35160
rect 23820 35040 24180 35160
rect 24300 35040 24420 35160
rect 24540 35040 24660 35160
rect 24780 35040 24900 35160
rect 25020 35040 25140 35160
rect 25260 35040 25620 35160
rect 25740 35040 25860 35160
rect 25980 35040 26100 35160
rect 26220 35040 26340 35160
rect 26460 35040 26820 35160
rect 26940 35040 27300 35160
rect 27420 35040 27540 35160
rect 27660 35040 27780 35160
rect 27900 35040 28020 35160
rect 28140 35040 28260 35160
rect 28380 35040 28500 35160
rect 28620 35040 28740 35160
rect 28860 35040 28980 35160
rect 29100 35040 29220 35160
rect 29340 35040 29460 35160
rect 29580 35040 29700 35160
rect 29820 35040 29940 35160
rect 30060 35040 30180 35160
rect 30300 35040 30420 35160
rect 30540 35040 30660 35160
rect 30780 35040 30900 35160
rect 31020 35040 31140 35160
rect 31260 35040 31620 35160
rect 31740 35040 31860 35160
rect 31980 35040 32340 35160
rect 32460 35040 32820 35160
rect 32940 35040 33060 35160
rect 33180 35040 33300 35160
rect 33420 35040 33540 35160
rect 33660 35040 33780 35160
rect 33900 35040 34020 35160
rect 34140 35040 34260 35160
rect 34380 35040 34500 35160
rect 34620 35040 34980 35160
rect 35100 35040 35220 35160
rect 35340 35040 35460 35160
rect 35580 35040 35700 35160
rect 35820 35040 35940 35160
rect 36060 35040 36180 35160
rect 36300 35040 36420 35160
rect 36540 35040 36660 35160
rect 36780 35040 36900 35160
rect 37020 35040 37140 35160
rect 37260 35040 37380 35160
rect 37500 35040 37620 35160
rect 37740 35040 37860 35160
rect 37980 35040 38100 35160
rect 38220 35040 38340 35160
rect 38460 35040 38580 35160
rect 38700 35040 38820 35160
rect 38940 35040 39300 35160
rect 39420 35040 39540 35160
rect 39660 35040 39780 35160
rect 39900 35040 40020 35160
rect 40140 35040 40500 35160
rect 40620 35040 40980 35160
rect 41100 35040 41220 35160
rect 41340 35040 41460 35160
rect 41580 35040 41940 35160
rect 42060 35040 42180 35160
rect 42300 35040 42420 35160
rect 42540 35040 42660 35160
rect 42780 35040 42900 35160
rect 43020 35040 43140 35160
rect 43260 35040 43380 35160
rect 43500 35040 43860 35160
rect 43980 35040 44100 35160
rect 44220 35040 44340 35160
rect 44460 35040 44580 35160
rect 44700 35040 44820 35160
rect 44940 35040 45060 35160
rect 45180 35040 45300 35160
rect 45420 35040 45540 35160
rect 45660 35040 45780 35160
rect 45900 35040 46020 35160
rect 46140 35040 46500 35160
rect 46620 35040 46740 35160
rect 46860 35040 46980 35160
rect 47100 35040 47220 35160
rect 47340 35040 47460 35160
rect 47580 35040 47700 35160
rect 47820 35040 47940 35160
rect 48060 35040 48180 35160
rect 48300 35040 48420 35160
rect 48540 35040 48660 35160
rect 48780 35040 48900 35160
rect 49020 35040 49140 35160
rect 49260 35040 49380 35160
rect 49500 35040 49620 35160
rect 49740 35040 49860 35160
rect 49980 35040 50100 35160
rect 50220 35040 53310 35160
rect 54180 35040 54240 35160
rect 1155 35010 54240 35040
rect 6630 34906 6750 35010
rect 6630 34320 6750 34334
rect 6870 34906 6990 34920
rect 6660 33810 6750 33990
rect 6540 33795 6750 33810
rect 5940 33720 6750 33795
rect 6840 33734 6870 33810
rect 6840 33720 6990 33734
rect 7260 34906 7380 35010
rect 7830 34906 7950 35010
rect 7830 34320 7950 34334
rect 8070 34906 8190 34920
rect 7860 33810 7950 33990
rect 7260 33720 7380 33734
rect 7740 33720 7950 33810
rect 8040 33734 8070 33810
rect 8040 33720 8190 33734
rect 8460 34906 8580 35010
rect 9210 34920 9330 35010
rect 8460 33720 8580 33734
rect 8940 34906 9060 34920
rect 9180 34860 9330 34920
rect 9180 33990 9194 34860
rect 9316 33990 9330 34860
rect 9180 33930 9330 33990
rect 9600 34906 9840 34920
rect 9060 33734 9150 33810
rect 8940 33720 9150 33734
rect 9600 33734 9660 34906
rect 9780 33810 9840 34906
rect 10110 34860 10260 35010
rect 11370 34920 11490 35010
rect 10110 33990 10124 34860
rect 10246 33990 10260 34860
rect 10110 33930 10260 33990
rect 10380 34906 10500 34920
rect 9780 33734 9900 33810
rect 9600 33720 9900 33734
rect 10260 33734 10380 33810
rect 10260 33720 10500 33734
rect 11100 34906 11220 34920
rect 11340 34860 11490 34920
rect 11340 33990 11354 34860
rect 11476 33990 11490 34860
rect 11340 33930 11490 33990
rect 11760 34906 12000 34920
rect 11220 33734 11310 33810
rect 11100 33720 11310 33734
rect 11760 33734 11820 34906
rect 11940 33810 12000 34906
rect 12270 34860 12420 35010
rect 12270 33990 12284 34860
rect 12406 33990 12420 34860
rect 12270 33930 12420 33990
rect 12540 34906 12660 34920
rect 11940 33734 12060 33810
rect 11760 33720 12060 33734
rect 12420 33734 12540 33810
rect 12420 33720 12660 33734
rect 13740 34890 13860 34920
rect 13980 34890 14100 35010
rect 15180 34906 15300 35010
rect 15180 34320 15300 34334
rect 15420 34906 15540 34920
rect 5940 33705 6660 33720
rect 6540 33690 6660 33705
rect 6840 33210 6930 33720
rect 7740 33690 7860 33720
rect 8040 33210 8130 33720
rect 9180 33630 9270 33720
rect 9180 33540 9570 33630
rect 9810 33510 9900 33720
rect 11340 33630 11430 33720
rect 11340 33540 11730 33630
rect 11970 33510 12060 33720
rect 9810 33420 10020 33510
rect 9360 33330 9630 33420
rect 9540 33240 9630 33330
rect 9750 33390 10020 33420
rect 9750 33330 9900 33390
rect 11970 33420 12180 33510
rect 11520 33330 11790 33420
rect 6660 33090 6930 33210
rect 7140 33150 7260 33180
rect 6570 32880 6660 33090
rect 7740 33195 8130 33210
rect 7620 33105 8130 33195
rect 8460 33195 8580 33210
rect 8460 33180 8700 33195
rect 7740 33090 8130 33105
rect 8340 33150 8700 33180
rect 6810 32880 7350 32940
rect 7770 32880 7860 33090
rect 8460 33105 8700 33150
rect 8460 33090 8580 33105
rect 8940 33090 9060 33210
rect 9180 33090 9450 33180
rect 9360 33030 9450 33090
rect 8010 32880 8550 32940
rect 8940 32880 9150 32970
rect 9360 32940 9420 33030
rect 6540 32866 6660 32880
rect 6540 32280 6660 32294
rect 6780 32866 7380 32880
rect 6900 32850 7260 32866
rect 6780 32280 6900 32294
rect 7020 32730 7140 32760
rect 7020 32190 7140 32310
rect 7260 32280 7380 32294
rect 7740 32866 7860 32880
rect 7740 32280 7860 32294
rect 7980 32866 8580 32880
rect 8100 32850 8460 32866
rect 7980 32280 8100 32294
rect 8220 32730 8340 32760
rect 8220 32190 8340 32310
rect 8460 32280 8580 32294
rect 8940 32866 9060 32880
rect 9750 32820 9840 33330
rect 11700 33240 11790 33330
rect 11910 33390 12180 33420
rect 11910 33330 12060 33390
rect 10380 33195 10500 33210
rect 10380 33105 10860 33195
rect 10380 33090 10500 33105
rect 11100 33090 11220 33210
rect 11340 33090 11610 33180
rect 9960 33030 10050 33090
rect 11520 33030 11610 33090
rect 10260 32880 10500 32970
rect 8940 32280 9060 32294
rect 9180 32746 9330 32790
rect 9180 32324 9194 32746
rect 9316 32324 9330 32746
rect 9180 32280 9330 32324
rect 9600 32760 9840 32820
rect 10380 32866 10500 32880
rect 9600 32340 9660 32760
rect 9780 32340 9840 32760
rect 9600 32280 9840 32340
rect 10110 32746 10260 32790
rect 10110 32324 10124 32746
rect 10246 32324 10260 32746
rect 9210 32190 9330 32280
rect 10110 32190 10260 32324
rect 10380 32280 10500 32294
rect 11100 32880 11310 32970
rect 11520 32940 11580 33030
rect 11100 32866 11220 32880
rect 11910 32820 12000 33330
rect 12540 33195 12660 33210
rect 13500 33195 13620 33210
rect 12540 33105 13620 33195
rect 12540 33090 12660 33105
rect 13500 33090 13620 33105
rect 12120 33030 12210 33090
rect 12420 32880 12660 32970
rect 11100 32280 11220 32294
rect 11340 32746 11490 32790
rect 11340 32324 11354 32746
rect 11476 32324 11490 32746
rect 11340 32280 11490 32324
rect 11760 32760 12000 32820
rect 12540 32866 12660 32880
rect 11760 32340 11820 32760
rect 11940 32340 12000 32760
rect 11760 32280 12000 32340
rect 12270 32746 12420 32790
rect 12270 32324 12284 32746
rect 12406 32324 12420 32746
rect 11370 32190 11490 32280
rect 12270 32190 12420 32324
rect 12540 32280 12660 32294
rect 13740 32550 13860 34320
rect 15420 34095 15540 34334
rect 15660 34906 15780 35010
rect 15660 34320 15780 34334
rect 16620 34906 16740 35010
rect 14100 34005 15540 34095
rect 13980 33195 14100 33210
rect 15180 33195 15300 33210
rect 13980 33105 15300 33195
rect 13980 33090 14100 33105
rect 15180 33090 15300 33105
rect 14100 32805 14940 32895
rect 15420 32880 15540 34005
rect 16620 33720 16740 33734
rect 17010 34906 17130 34920
rect 17250 34906 17370 35010
rect 17250 34320 17370 34334
rect 19260 34906 19380 35010
rect 19260 34320 19380 34334
rect 19500 34906 19620 34920
rect 17250 33810 17340 33990
rect 17130 33734 17160 33810
rect 17010 33720 17160 33734
rect 17250 33795 17460 33810
rect 17250 33720 18300 33795
rect 16860 33390 16980 33510
rect 17070 33210 17160 33720
rect 17340 33705 18300 33720
rect 17340 33690 17460 33705
rect 18540 33795 18660 33810
rect 19260 33795 19380 33810
rect 18540 33705 19380 33795
rect 18540 33690 18660 33705
rect 19260 33690 19380 33705
rect 16620 33195 16740 33210
rect 16500 33180 16740 33195
rect 16500 33150 16860 33180
rect 16500 33105 16740 33150
rect 16620 33090 16740 33105
rect 17070 33090 17460 33210
rect 16650 32880 17190 32940
rect 17340 32880 17430 33090
rect 19500 32880 19620 34334
rect 19740 34906 19860 35010
rect 19740 34320 19860 34334
rect 20700 34906 20820 34920
rect 20700 34320 20820 34334
rect 20940 34906 21060 35010
rect 20940 34320 21060 34334
rect 21180 34906 21300 34920
rect 21180 34320 21300 34334
rect 21420 34906 21540 35010
rect 21420 34320 21540 34334
rect 23340 34906 23460 35010
rect 20700 34110 20790 34320
rect 21180 34230 21270 34320
rect 20910 34140 21270 34230
rect 19740 34095 19860 34110
rect 20700 34095 20820 34110
rect 19740 34005 20820 34095
rect 19740 33990 19860 34005
rect 20700 33990 20820 34005
rect 19740 33195 19860 33210
rect 19740 33105 19980 33195
rect 19740 33090 19860 33105
rect 15180 32866 15300 32880
rect 13980 32550 14100 32580
rect 13980 32190 14100 32280
rect 15420 32866 15690 32880
rect 15420 32790 15570 32866
rect 15180 32190 15300 32294
rect 15570 32280 15690 32294
rect 16620 32866 17220 32880
rect 16740 32850 17100 32866
rect 16620 32280 16740 32294
rect 16860 32730 16980 32760
rect 16860 32190 16980 32310
rect 17100 32280 17220 32294
rect 17340 32866 17460 32880
rect 17340 32280 17460 32294
rect 19350 32866 19620 32880
rect 19470 32790 19620 32866
rect 19740 32866 19860 32880
rect 19350 32280 19470 32294
rect 20700 32670 20790 33990
rect 20910 33090 21000 34140
rect 21090 33690 21300 33810
rect 23340 33720 23460 33734
rect 23730 34906 23850 34920
rect 23970 34906 24090 35010
rect 23970 34320 24090 34334
rect 24780 34906 24900 35010
rect 23970 33810 24060 33990
rect 23850 33734 23880 33810
rect 23730 33720 23880 33734
rect 23970 33795 24180 33810
rect 24540 33795 24660 33810
rect 23970 33720 24660 33795
rect 24780 33720 24900 33734
rect 25170 34906 25290 34920
rect 25410 34906 25530 35010
rect 26250 34920 26370 35010
rect 25410 34320 25530 34334
rect 25980 34906 26100 34920
rect 25290 33734 25320 33810
rect 25170 33720 25320 33734
rect 25410 33720 25500 33990
rect 22395 33405 22860 33495
rect 21420 33195 21540 33210
rect 22395 33195 22485 33405
rect 22980 33405 23340 33495
rect 23790 33210 23880 33720
rect 24060 33705 24660 33720
rect 24060 33690 24180 33705
rect 24540 33690 24660 33705
rect 25020 33495 25140 33510
rect 24180 33405 25140 33495
rect 25020 33390 25140 33405
rect 25230 33210 25320 33720
rect 26220 34860 26370 34920
rect 26220 33990 26234 34860
rect 26356 33990 26370 34860
rect 26220 33930 26370 33990
rect 26640 34906 26880 34920
rect 26100 33734 26250 33810
rect 25980 33720 26250 33734
rect 26640 33734 26700 34906
rect 26820 33734 26880 34906
rect 27150 34860 27300 35010
rect 27150 33990 27164 34860
rect 27286 33990 27300 34860
rect 27150 33930 27300 33990
rect 27420 34906 27540 34920
rect 26640 33720 26880 33734
rect 27300 33734 27420 33810
rect 27300 33720 27540 33734
rect 30300 34890 30420 34920
rect 30540 34890 30660 35010
rect 31020 34906 31140 35010
rect 31020 34320 31140 34334
rect 31260 34906 31380 34920
rect 26730 33510 26820 33720
rect 26700 33390 26820 33510
rect 21420 33105 22485 33195
rect 21420 33090 21540 33105
rect 23340 33195 23460 33210
rect 22740 33180 23460 33195
rect 22740 33150 23580 33180
rect 22740 33105 23460 33150
rect 23340 33090 23460 33105
rect 21000 33000 21330 33090
rect 23790 33090 24180 33210
rect 24780 33195 24900 33210
rect 24420 33180 24900 33195
rect 24420 33150 25020 33180
rect 24420 33105 24900 33150
rect 24780 33090 24900 33105
rect 21240 32970 21330 33000
rect 21240 32880 21510 32970
rect 23370 32880 23910 32940
rect 24060 32880 24150 33090
rect 25230 33090 25260 33210
rect 25380 33090 25620 33210
rect 25740 33195 25860 33210
rect 25980 33195 26100 33210
rect 25740 33105 26100 33195
rect 25740 33090 25860 33105
rect 25980 33090 26100 33105
rect 26220 33150 26520 33240
rect 26730 33210 26820 33390
rect 26220 33120 26310 33150
rect 26730 33120 26880 33210
rect 24810 32880 25350 32940
rect 25500 32880 25590 33090
rect 25980 32880 26250 32970
rect 21030 32866 21150 32880
rect 20700 32580 20910 32670
rect 19740 32190 19860 32294
rect 20790 32566 20910 32580
rect 20790 32280 20910 32294
rect 21030 32190 21150 32294
rect 21420 32866 21540 32880
rect 21420 32280 21540 32294
rect 23340 32866 23940 32880
rect 23460 32850 23820 32866
rect 23340 32280 23460 32294
rect 23580 32730 23700 32760
rect 23580 32190 23700 32310
rect 23820 32280 23940 32294
rect 24060 32866 24180 32880
rect 24060 32280 24180 32294
rect 24780 32866 25380 32880
rect 24900 32850 25260 32866
rect 24780 32280 24900 32294
rect 25020 32730 25140 32760
rect 25020 32190 25140 32310
rect 25260 32280 25380 32294
rect 25500 32866 25620 32880
rect 25500 32280 25620 32294
rect 25980 32866 26100 32880
rect 26790 32820 26880 33120
rect 27000 33030 27090 33090
rect 27300 32880 27540 32970
rect 25980 32280 26100 32294
rect 26220 32746 26370 32790
rect 26220 32324 26234 32746
rect 26356 32324 26370 32746
rect 26220 32280 26370 32324
rect 26640 32760 26880 32820
rect 27420 32866 27540 32880
rect 26640 32340 26700 32760
rect 26820 32340 26880 32760
rect 26640 32280 26880 32340
rect 27150 32746 27300 32790
rect 27150 32324 27164 32746
rect 27286 32324 27300 32746
rect 26250 32190 26370 32280
rect 27150 32190 27300 32324
rect 27420 32280 27540 32294
rect 30300 32550 30420 34320
rect 31260 33795 31380 34334
rect 31500 34906 31620 35010
rect 31500 34320 31620 34334
rect 31980 34906 32100 35010
rect 31740 33795 31860 33810
rect 31260 33705 31860 33795
rect 31980 33720 32100 33734
rect 32370 34906 32490 34920
rect 32610 34906 32730 35010
rect 32610 34320 32730 34334
rect 33180 34906 33300 35010
rect 33180 34320 33300 34334
rect 33420 34906 33540 34920
rect 32610 33810 32700 33990
rect 32490 33734 32520 33810
rect 32370 33720 32520 33734
rect 32610 33720 32820 33810
rect 31260 32880 31380 33705
rect 31740 33690 31860 33705
rect 31620 33405 31980 33495
rect 32220 33495 32340 33510
rect 32100 33405 32340 33495
rect 32220 33390 32340 33405
rect 32430 33210 32520 33720
rect 32700 33690 32820 33720
rect 31980 33195 32100 33210
rect 31860 33180 32100 33195
rect 32430 33195 32820 33210
rect 31860 33150 32220 33180
rect 31860 33105 32100 33150
rect 31980 33090 32100 33105
rect 32430 33105 32940 33195
rect 32430 33090 32820 33105
rect 33180 33090 33300 33210
rect 32010 32880 32550 32940
rect 32700 32880 32790 33090
rect 33420 32880 33540 34334
rect 33660 34906 33780 35010
rect 33660 34320 33780 34334
rect 34620 34906 34740 35010
rect 34620 34320 34740 34334
rect 34860 34906 34980 34920
rect 33660 33690 33780 33810
rect 34860 32880 34980 34334
rect 35100 34906 35220 35010
rect 35100 34320 35220 34334
rect 36060 34906 36180 35010
rect 36060 34320 36180 34334
rect 36300 34906 36420 34920
rect 36060 33195 36180 33210
rect 35460 33105 36180 33195
rect 36060 33090 36180 33105
rect 36300 32880 36420 34334
rect 36540 34906 36660 35010
rect 36540 34320 36660 34334
rect 37500 34906 37620 35010
rect 37500 34320 37620 34334
rect 37740 34906 37860 34920
rect 37740 34095 37860 34334
rect 37980 34906 38100 35010
rect 37980 34320 38100 34334
rect 38940 34906 39060 35010
rect 38940 34320 39060 34334
rect 39180 34906 39300 34920
rect 37740 34005 38700 34095
rect 36540 33795 36660 33810
rect 37500 33795 37620 33810
rect 36540 33705 37620 33795
rect 36540 33690 36660 33705
rect 37500 33690 37620 33705
rect 37740 32880 37860 34005
rect 38940 33195 39060 33210
rect 38340 33105 39060 33195
rect 38940 33090 39060 33105
rect 39180 32895 39300 34334
rect 39420 34906 39540 35010
rect 39420 34320 39540 34334
rect 40140 34906 40260 35010
rect 40140 33720 40260 33734
rect 40530 34906 40650 34920
rect 40770 34906 40890 35010
rect 40770 34320 40890 34334
rect 41580 34906 41700 35010
rect 41580 34320 41700 34334
rect 41820 34906 41940 34920
rect 40770 33810 40860 33990
rect 40650 33734 40680 33810
rect 40530 33720 40680 33734
rect 40770 33795 40980 33810
rect 40770 33720 41580 33795
rect 40590 33210 40680 33720
rect 40860 33705 41580 33720
rect 40860 33690 40980 33705
rect 39420 33195 39540 33210
rect 40140 33195 40260 33210
rect 39420 33180 40260 33195
rect 39420 33150 40380 33180
rect 39420 33105 40260 33150
rect 39420 33090 39540 33105
rect 40140 33090 40260 33105
rect 40590 33090 40980 33210
rect 41580 33195 41700 33210
rect 41460 33105 41700 33195
rect 41580 33090 41700 33105
rect 39900 32895 40020 32910
rect 31110 32866 31380 32880
rect 30540 32550 30660 32580
rect 31230 32790 31380 32866
rect 31500 32866 31620 32880
rect 31110 32280 31230 32294
rect 30540 32190 30660 32280
rect 31500 32190 31620 32294
rect 31980 32866 32580 32880
rect 32100 32850 32460 32866
rect 31980 32280 32100 32294
rect 32220 32730 32340 32760
rect 32220 32190 32340 32310
rect 32460 32280 32580 32294
rect 32700 32866 32820 32880
rect 32700 32280 32820 32294
rect 33180 32866 33300 32880
rect 33420 32866 33690 32880
rect 33420 32790 33570 32866
rect 33180 32190 33300 32294
rect 33570 32280 33690 32294
rect 34620 32866 34740 32880
rect 34860 32866 35130 32880
rect 34860 32790 35010 32866
rect 34620 32190 34740 32294
rect 35010 32280 35130 32294
rect 36060 32866 36180 32880
rect 36300 32866 36570 32880
rect 36300 32790 36450 32866
rect 36060 32190 36180 32294
rect 36450 32280 36570 32294
rect 37590 32866 37860 32880
rect 37710 32790 37860 32866
rect 37980 32866 38100 32880
rect 37590 32280 37710 32294
rect 37980 32190 38100 32294
rect 38940 32866 39060 32880
rect 39180 32866 40020 32895
rect 40170 32880 40710 32940
rect 40860 32880 40950 33090
rect 41820 32880 41940 34334
rect 42060 34906 42180 35010
rect 42060 34320 42180 34334
rect 43020 34906 43140 35010
rect 43020 33720 43140 33734
rect 43410 34906 43530 34920
rect 43650 34906 43770 35010
rect 44490 34920 44610 35010
rect 43650 34320 43770 34334
rect 44220 34906 44340 34920
rect 43650 33810 43740 33990
rect 43530 33734 43560 33810
rect 43410 33720 43560 33734
rect 43650 33720 43860 33810
rect 44460 34860 44610 34920
rect 44460 33990 44474 34860
rect 44596 33990 44610 34860
rect 44460 33930 44610 33990
rect 44880 34906 45120 34920
rect 44340 33734 44490 33810
rect 44220 33720 44490 33734
rect 44880 33734 44940 34906
rect 45060 33734 45120 34906
rect 45390 34860 45540 35010
rect 45390 33990 45404 34860
rect 45526 33990 45540 34860
rect 45390 33930 45540 33990
rect 45660 34906 45780 34920
rect 44880 33720 45120 33734
rect 45540 33734 45660 33810
rect 45540 33720 45780 33734
rect 46140 34906 46260 35010
rect 46140 33720 46260 33734
rect 46530 34906 46650 34920
rect 46770 34906 46890 35010
rect 46770 34320 46890 34334
rect 47580 34906 47700 35010
rect 47580 34320 47700 34334
rect 47820 34906 47940 34920
rect 46770 33810 46860 33990
rect 46650 33734 46680 33810
rect 46530 33720 46680 33734
rect 46770 33795 46980 33810
rect 47340 33795 47460 33810
rect 46770 33720 47460 33795
rect 42300 33495 42420 33510
rect 43260 33495 43380 33510
rect 42300 33405 43380 33495
rect 42300 33390 42420 33405
rect 43260 33390 43380 33405
rect 43470 33210 43560 33720
rect 43740 33690 43860 33720
rect 44970 33510 45060 33720
rect 44940 33390 45060 33510
rect 46380 33495 46500 33510
rect 46020 33405 46500 33495
rect 46380 33390 46500 33405
rect 42060 33195 42180 33210
rect 43020 33195 43140 33210
rect 42060 33180 43140 33195
rect 42060 33150 43260 33180
rect 42060 33105 43140 33150
rect 42060 33090 42180 33105
rect 43020 33090 43140 33105
rect 43470 33090 43500 33210
rect 43620 33090 43860 33210
rect 43980 33195 44100 33210
rect 44220 33195 44340 33210
rect 43980 33105 44340 33195
rect 43980 33090 44100 33105
rect 44220 33090 44340 33105
rect 44460 33150 44760 33240
rect 44970 33210 45060 33390
rect 46590 33210 46680 33720
rect 46860 33705 47460 33720
rect 46860 33690 46980 33705
rect 47340 33690 47460 33705
rect 47820 33795 47940 34334
rect 48060 34906 48180 35010
rect 48060 34320 48180 34334
rect 49020 34906 49140 35010
rect 49020 34320 49140 34334
rect 49260 34906 49380 34920
rect 49020 33795 49140 33810
rect 47820 33705 49140 33795
rect 44460 33120 44550 33150
rect 44970 33120 45120 33210
rect 43050 32880 43590 32940
rect 43740 32880 43830 33090
rect 44220 32880 44490 32970
rect 39180 32790 39330 32866
rect 38940 32190 39060 32294
rect 39450 32805 40020 32866
rect 39900 32790 40020 32805
rect 40140 32866 40740 32880
rect 39330 32280 39450 32294
rect 40260 32850 40620 32866
rect 40140 32280 40260 32294
rect 40380 32730 40500 32760
rect 40380 32190 40500 32310
rect 40620 32280 40740 32294
rect 40860 32866 40980 32880
rect 41580 32866 41700 32880
rect 41340 32595 41460 32610
rect 40980 32505 41460 32595
rect 41340 32490 41460 32505
rect 40860 32280 40980 32294
rect 41820 32866 42090 32880
rect 41820 32790 41970 32866
rect 41580 32190 41700 32294
rect 41970 32280 42090 32294
rect 43020 32866 43620 32880
rect 43140 32850 43500 32866
rect 43020 32280 43140 32294
rect 43260 32730 43380 32760
rect 43260 32190 43380 32310
rect 43500 32280 43620 32294
rect 43740 32866 43860 32880
rect 43740 32280 43860 32294
rect 44220 32866 44340 32880
rect 45030 32820 45120 33120
rect 46260 33150 46380 33180
rect 45240 33030 45330 33090
rect 46590 33090 46980 33210
rect 45540 32880 45780 32970
rect 46170 32880 46710 32940
rect 46860 32880 46950 33090
rect 47820 32880 47940 33705
rect 49020 33690 49140 33705
rect 49260 33495 49380 34334
rect 49500 34906 49620 35010
rect 49500 34320 49620 34334
rect 48180 33405 49380 33495
rect 48180 33105 48300 33195
rect 49260 32880 49380 33405
rect 44220 32280 44340 32294
rect 44460 32746 44610 32790
rect 44460 32324 44474 32746
rect 44596 32324 44610 32746
rect 44460 32280 44610 32324
rect 44880 32760 45120 32820
rect 45660 32866 45780 32880
rect 44880 32340 44940 32760
rect 45060 32340 45120 32760
rect 44880 32280 45120 32340
rect 45390 32746 45540 32790
rect 45390 32324 45404 32746
rect 45526 32324 45540 32746
rect 44490 32190 44610 32280
rect 45390 32190 45540 32324
rect 45660 32280 45780 32294
rect 46140 32866 46740 32880
rect 46260 32850 46620 32866
rect 46140 32280 46260 32294
rect 46380 32730 46500 32760
rect 46380 32190 46500 32310
rect 46620 32280 46740 32294
rect 46860 32866 46980 32880
rect 46860 32280 46980 32294
rect 47670 32866 47940 32880
rect 47790 32790 47940 32866
rect 48060 32866 48180 32880
rect 47670 32280 47790 32294
rect 48060 32190 48180 32294
rect 49110 32866 49380 32880
rect 49230 32790 49380 32866
rect 49500 32866 49620 32880
rect 49110 32280 49230 32294
rect 49500 32190 49620 32294
rect 3135 32160 52260 32190
rect 3135 32040 3194 32160
rect 4066 32040 5220 32160
rect 5340 32040 5460 32160
rect 5580 32040 5700 32160
rect 5820 32040 5940 32160
rect 6060 32040 6180 32160
rect 6300 32040 6420 32160
rect 6540 32040 6900 32160
rect 7020 32040 7140 32160
rect 7260 32040 7380 32160
rect 7500 32040 7620 32160
rect 7740 32040 7860 32160
rect 7980 32040 8100 32160
rect 8220 32040 8340 32160
rect 8460 32040 8580 32160
rect 8700 32040 8820 32160
rect 8940 32040 9060 32160
rect 9180 32040 9300 32160
rect 9420 32040 9540 32160
rect 9660 32040 9780 32160
rect 9900 32040 10260 32160
rect 10380 32040 10500 32160
rect 10620 32040 10740 32160
rect 10860 32040 10980 32160
rect 11100 32040 11460 32160
rect 11580 32040 11940 32160
rect 12060 32040 12420 32160
rect 12540 32040 12660 32160
rect 12780 32040 12900 32160
rect 13020 32040 13140 32160
rect 13260 32040 13380 32160
rect 13500 32040 13620 32160
rect 13740 32040 13860 32160
rect 13980 32040 14100 32160
rect 14220 32040 14340 32160
rect 14460 32040 14580 32160
rect 14700 32040 14820 32160
rect 14940 32040 15060 32160
rect 15180 32040 15540 32160
rect 15660 32040 15780 32160
rect 15900 32040 16020 32160
rect 16140 32040 16260 32160
rect 16380 32040 16500 32160
rect 16620 32040 16740 32160
rect 16860 32040 16980 32160
rect 17100 32040 17460 32160
rect 17580 32040 17700 32160
rect 17820 32040 17940 32160
rect 18060 32040 18180 32160
rect 18300 32040 18420 32160
rect 18540 32040 18660 32160
rect 18780 32040 18900 32160
rect 19020 32040 19140 32160
rect 19260 32040 19380 32160
rect 19500 32040 19620 32160
rect 19740 32040 19860 32160
rect 19980 32040 20100 32160
rect 20220 32040 20340 32160
rect 20460 32040 20580 32160
rect 20700 32040 20820 32160
rect 20940 32040 21060 32160
rect 21180 32040 21540 32160
rect 21660 32040 21780 32160
rect 21900 32040 22020 32160
rect 22140 32040 22260 32160
rect 22380 32040 22500 32160
rect 22620 32040 22740 32160
rect 22860 32040 22980 32160
rect 23100 32040 23220 32160
rect 23340 32040 23460 32160
rect 23580 32040 23700 32160
rect 23820 32040 24180 32160
rect 24300 32040 24420 32160
rect 24540 32040 24660 32160
rect 24780 32040 25140 32160
rect 25260 32040 25620 32160
rect 25740 32040 25860 32160
rect 25980 32040 26340 32160
rect 26460 32040 26820 32160
rect 26940 32040 27060 32160
rect 27180 32040 27300 32160
rect 27420 32040 27540 32160
rect 27660 32040 27780 32160
rect 27900 32040 28020 32160
rect 28140 32040 28260 32160
rect 28380 32040 28500 32160
rect 28620 32040 28740 32160
rect 28860 32040 28980 32160
rect 29100 32040 29220 32160
rect 29340 32040 29460 32160
rect 29580 32040 29700 32160
rect 29820 32040 29940 32160
rect 30060 32040 30180 32160
rect 30300 32040 30420 32160
rect 30540 32040 30660 32160
rect 30780 32040 30900 32160
rect 31020 32040 31140 32160
rect 31260 32040 31380 32160
rect 31500 32040 31620 32160
rect 31740 32040 31860 32160
rect 31980 32040 32340 32160
rect 32460 32040 32580 32160
rect 32700 32040 32820 32160
rect 32940 32040 33060 32160
rect 33180 32040 33540 32160
rect 33660 32040 33780 32160
rect 33900 32040 34020 32160
rect 34140 32040 34260 32160
rect 34380 32040 34500 32160
rect 34620 32040 34980 32160
rect 35100 32040 35220 32160
rect 35340 32040 35460 32160
rect 35580 32040 35700 32160
rect 35820 32040 35940 32160
rect 36060 32040 36420 32160
rect 36540 32040 36660 32160
rect 36780 32040 36900 32160
rect 37020 32040 37140 32160
rect 37260 32040 37380 32160
rect 37500 32040 37620 32160
rect 37740 32040 38100 32160
rect 38220 32040 38340 32160
rect 38460 32040 38580 32160
rect 38700 32040 38820 32160
rect 38940 32040 39300 32160
rect 39420 32040 39540 32160
rect 39660 32040 39780 32160
rect 39900 32040 40020 32160
rect 40140 32040 40260 32160
rect 40380 32040 40500 32160
rect 40620 32040 40980 32160
rect 41100 32040 41220 32160
rect 41340 32040 41460 32160
rect 41580 32040 41700 32160
rect 41820 32040 41940 32160
rect 42060 32040 42180 32160
rect 42300 32040 42420 32160
rect 42540 32040 42660 32160
rect 42780 32040 42900 32160
rect 43020 32040 43380 32160
rect 43500 32040 43860 32160
rect 43980 32040 44100 32160
rect 44220 32040 44340 32160
rect 44460 32040 44580 32160
rect 44700 32040 44820 32160
rect 44940 32040 45060 32160
rect 45180 32040 45300 32160
rect 45420 32040 45540 32160
rect 45660 32040 45780 32160
rect 45900 32040 46020 32160
rect 46140 32040 46260 32160
rect 46380 32040 46500 32160
rect 46620 32040 46740 32160
rect 46860 32040 46980 32160
rect 47100 32040 47220 32160
rect 47340 32040 47460 32160
rect 47580 32040 47700 32160
rect 47820 32040 47940 32160
rect 48060 32040 48180 32160
rect 48300 32040 48420 32160
rect 48540 32040 48660 32160
rect 48780 32040 48900 32160
rect 49020 32040 49140 32160
rect 49260 32040 49380 32160
rect 49500 32040 49620 32160
rect 49740 32040 49860 32160
rect 49980 32040 50100 32160
rect 50220 32040 51330 32160
rect 52200 32040 52260 32160
rect 3135 32010 52260 32040
rect 5340 31906 5460 31920
rect 5580 31876 5730 32010
rect 6510 31920 6630 32010
rect 5580 31454 5594 31876
rect 5716 31454 5730 31876
rect 5580 31410 5730 31454
rect 6000 31860 6240 31920
rect 6000 31440 6060 31860
rect 6180 31440 6240 31860
rect 5340 31320 5460 31334
rect 6000 31380 6240 31440
rect 6510 31876 6660 31920
rect 6510 31454 6524 31876
rect 6646 31454 6660 31876
rect 6510 31410 6660 31454
rect 6780 31906 6900 31920
rect 5340 31230 5580 31320
rect 5790 31110 5880 31170
rect 6000 30870 6090 31380
rect 6780 31320 6900 31334
rect 7980 31906 8100 31920
rect 8220 31890 8340 32010
rect 8220 31440 8340 31470
rect 8460 31906 8580 31920
rect 8100 31334 8460 31350
rect 7980 31320 8580 31334
rect 8700 31906 8820 31920
rect 8700 31320 8820 31334
rect 9750 31906 9870 31920
rect 10140 31906 10260 32010
rect 11370 31920 11490 32010
rect 9870 31334 10020 31410
rect 9750 31320 10020 31334
rect 10140 31320 10260 31334
rect 11100 31906 11220 31920
rect 11340 31876 11490 31920
rect 11340 31454 11354 31876
rect 11476 31454 11490 31876
rect 11340 31410 11490 31454
rect 11760 31860 12000 31920
rect 11760 31440 11820 31860
rect 11940 31440 12000 31860
rect 11760 31380 12000 31440
rect 12270 31876 12420 32010
rect 14970 31920 15090 32010
rect 12270 31454 12284 31876
rect 12406 31454 12420 31876
rect 12270 31410 12420 31454
rect 12540 31906 12660 31920
rect 11100 31320 11220 31334
rect 6420 31170 6480 31260
rect 6690 31230 6900 31320
rect 8010 31260 8550 31320
rect 6390 31110 6480 31170
rect 6390 31020 6660 31110
rect 6780 30990 6900 31110
rect 7980 31095 8100 31110
rect 7140 31050 8100 31095
rect 8700 31110 8790 31320
rect 7140 31020 8220 31050
rect 7140 31005 8100 31020
rect 7980 30990 8100 31005
rect 8430 30990 8460 31110
rect 8580 30990 8820 31110
rect 5940 30810 6090 30870
rect 5820 30780 6090 30810
rect 6210 30870 6300 30960
rect 6210 30780 6480 30870
rect 5820 30690 6030 30780
rect 8220 30690 8340 30810
rect 5940 30480 6030 30690
rect 6270 30570 6660 30660
rect 6570 30480 6660 30570
rect 8430 30480 8520 30990
rect 8700 30495 8820 30510
rect 8700 30480 8940 30495
rect 5340 30466 5580 30480
rect 5460 30390 5580 30466
rect 5940 30466 6240 30480
rect 5940 30390 6060 30466
rect 5340 29280 5460 29294
rect 5580 30210 5730 30270
rect 5580 29340 5594 30210
rect 5716 29340 5730 30210
rect 5580 29190 5730 29340
rect 6000 29294 6060 30390
rect 6180 29294 6240 30466
rect 6690 30466 6900 30480
rect 6690 30390 6780 30466
rect 6000 29280 6240 29294
rect 6510 30210 6660 30270
rect 6510 29340 6524 30210
rect 6646 29340 6660 30210
rect 6510 29280 6660 29340
rect 6780 29280 6900 29294
rect 7980 30466 8100 30480
rect 6510 29190 6630 29280
rect 7980 29190 8100 29294
rect 8370 30466 8520 30480
rect 8490 30390 8520 30466
rect 8610 30405 8940 30480
rect 8610 30390 8820 30405
rect 9660 30495 9780 30510
rect 9300 30405 9780 30495
rect 9660 30390 9780 30405
rect 8610 30210 8700 30390
rect 8370 29280 8490 29294
rect 8610 29866 8730 29880
rect 8610 29190 8730 29294
rect 9660 29866 9780 29880
rect 9660 29190 9780 29294
rect 9900 29866 10020 31320
rect 11100 31230 11370 31320
rect 11910 31080 12000 31380
rect 12540 31320 12660 31334
rect 12420 31230 12660 31320
rect 14700 31906 14820 31920
rect 14940 31876 15090 31920
rect 14940 31454 14954 31876
rect 15076 31454 15090 31876
rect 14940 31410 15090 31454
rect 15360 31860 15600 31920
rect 15360 31440 15420 31860
rect 15540 31440 15600 31860
rect 15360 31380 15600 31440
rect 15870 31876 16020 32010
rect 17370 31920 17490 32010
rect 15870 31454 15884 31876
rect 16006 31454 16020 31876
rect 15870 31410 16020 31454
rect 16140 31906 16260 31920
rect 14700 31320 14820 31334
rect 14700 31230 14910 31320
rect 11340 31050 11430 31080
rect 11340 30960 11640 31050
rect 11850 30990 12000 31080
rect 12120 31110 12210 31170
rect 15120 31170 15180 31260
rect 15120 31110 15210 31170
rect 12540 31095 12660 31110
rect 12540 31005 12780 31095
rect 12540 30990 12660 31005
rect 14700 31095 14820 31110
rect 14100 31005 14820 31095
rect 14700 30990 14820 31005
rect 14940 31020 15210 31110
rect 11850 30810 11940 30990
rect 15300 30870 15390 30960
rect 11820 30690 11940 30810
rect 15120 30780 15390 30870
rect 15510 30870 15600 31380
rect 16140 31320 16260 31334
rect 16020 31230 16260 31320
rect 17100 31906 17220 31920
rect 17340 31876 17490 31920
rect 17340 31454 17354 31876
rect 17476 31454 17490 31876
rect 17340 31410 17490 31454
rect 17760 31860 18000 31920
rect 17760 31440 17820 31860
rect 17940 31440 18000 31860
rect 17760 31380 18000 31440
rect 18270 31876 18420 32010
rect 19530 31920 19650 32010
rect 18270 31454 18284 31876
rect 18406 31454 18420 31876
rect 18270 31410 18420 31454
rect 18540 31906 18660 31920
rect 17100 31320 17220 31334
rect 17100 31230 17310 31320
rect 15720 31110 15810 31170
rect 17520 31170 17580 31260
rect 17520 31110 17610 31170
rect 16140 31095 16260 31110
rect 16140 31005 16860 31095
rect 16140 30990 16260 31005
rect 17340 31020 17610 31110
rect 17700 30870 17790 30960
rect 15510 30810 15660 30870
rect 15510 30780 15780 30810
rect 15570 30690 15780 30780
rect 17520 30780 17790 30870
rect 17910 30870 18000 31380
rect 18540 31320 18660 31334
rect 18420 31230 18660 31320
rect 19260 31906 19380 31920
rect 19500 31876 19650 31920
rect 19500 31454 19514 31876
rect 19636 31454 19650 31876
rect 19500 31410 19650 31454
rect 19920 31860 20160 31920
rect 19920 31440 19980 31860
rect 20100 31440 20160 31860
rect 19920 31380 20160 31440
rect 20430 31876 20580 32010
rect 20430 31454 20444 31876
rect 20566 31454 20580 31876
rect 20430 31410 20580 31454
rect 20700 31906 20820 31920
rect 19260 31320 19380 31334
rect 19260 31230 19530 31320
rect 18120 31110 18210 31170
rect 18540 31095 18660 31110
rect 18540 31005 19020 31095
rect 18540 30990 18660 31005
rect 20070 31080 20160 31380
rect 20700 31320 20820 31334
rect 21180 31906 21300 32010
rect 21570 31906 21690 31920
rect 21180 31320 21300 31334
rect 21420 31334 21570 31410
rect 21420 31320 21690 31334
rect 22140 31906 22260 31920
rect 22140 31320 22260 31334
rect 22380 31906 22500 31920
rect 22620 31890 22740 32010
rect 24060 31920 24180 32010
rect 22620 31440 22740 31470
rect 22860 31906 22980 31920
rect 22500 31334 22860 31350
rect 23700 31650 23820 31695
rect 23700 31605 23940 31650
rect 24060 31620 24180 31650
rect 24870 31906 24990 31920
rect 24870 31620 24990 31634
rect 22380 31320 22980 31334
rect 20580 31230 20820 31320
rect 19500 31050 19590 31080
rect 19500 30960 19800 31050
rect 20010 30990 20160 31080
rect 20280 31110 20370 31170
rect 20700 31095 20820 31110
rect 20940 31095 21060 31110
rect 20700 31005 21060 31095
rect 20700 30990 20820 31005
rect 20940 30990 21060 31005
rect 17910 30810 18060 30870
rect 20010 30810 20100 30990
rect 17910 30780 18180 30810
rect 17970 30690 18180 30780
rect 11850 30480 11940 30690
rect 14940 30570 15330 30660
rect 14940 30480 15030 30570
rect 15570 30480 15660 30690
rect 17340 30570 17730 30660
rect 17340 30480 17430 30570
rect 17970 30480 18060 30690
rect 19980 30690 20100 30810
rect 20010 30480 20100 30690
rect 11100 30466 11370 30480
rect 9900 29280 10020 29294
rect 10140 29866 10260 29880
rect 10140 29190 10260 29294
rect 11220 30390 11370 30466
rect 11760 30466 12000 30480
rect 11100 29280 11220 29294
rect 11340 30210 11490 30270
rect 11340 29340 11354 30210
rect 11476 29340 11490 30210
rect 11340 29280 11490 29340
rect 11760 29294 11820 30466
rect 11940 29294 12000 30466
rect 12420 30466 12660 30480
rect 12420 30390 12540 30466
rect 11760 29280 12000 29294
rect 12270 30210 12420 30270
rect 12270 29340 12284 30210
rect 12406 29340 12420 30210
rect 11370 29190 11490 29280
rect 12270 29190 12420 29340
rect 12540 29280 12660 29294
rect 14700 30466 14910 30480
rect 14820 30390 14910 30466
rect 15360 30466 15660 30480
rect 14700 29280 14820 29294
rect 14940 30210 15090 30270
rect 14940 29340 14954 30210
rect 15076 29340 15090 30210
rect 14940 29280 15090 29340
rect 15360 29294 15420 30466
rect 15540 30390 15660 30466
rect 15540 29294 15600 30390
rect 16020 30466 16260 30480
rect 16020 30390 16140 30466
rect 15360 29280 15600 29294
rect 15870 30210 16020 30270
rect 15870 29340 15884 30210
rect 16006 29340 16020 30210
rect 14970 29190 15090 29280
rect 15870 29190 16020 29340
rect 16140 29280 16260 29294
rect 17100 30466 17310 30480
rect 17220 30390 17310 30466
rect 17760 30466 18060 30480
rect 17100 29280 17220 29294
rect 17340 30210 17490 30270
rect 17340 29340 17354 30210
rect 17476 29340 17490 30210
rect 17340 29280 17490 29340
rect 17760 29294 17820 30466
rect 17940 30390 18060 30466
rect 17940 29294 18000 30390
rect 18420 30466 18660 30480
rect 18420 30390 18540 30466
rect 17760 29280 18000 29294
rect 18270 30210 18420 30270
rect 18270 29340 18284 30210
rect 18406 29340 18420 30210
rect 17370 29190 17490 29280
rect 18270 29190 18420 29340
rect 18540 29280 18660 29294
rect 19260 30466 19530 30480
rect 19380 30390 19530 30466
rect 19920 30466 20160 30480
rect 19260 29280 19380 29294
rect 19500 30210 19650 30270
rect 19500 29340 19514 30210
rect 19636 29340 19650 30210
rect 19500 29280 19650 29340
rect 19920 29294 19980 30466
rect 20100 29294 20160 30466
rect 20580 30466 20820 30480
rect 20580 30390 20700 30466
rect 19920 29280 20160 29294
rect 20430 30210 20580 30270
rect 20430 29340 20444 30210
rect 20566 29340 20580 30210
rect 19530 29190 19650 29280
rect 20430 29190 20580 29340
rect 20700 29280 20820 29294
rect 21180 29866 21300 29880
rect 21180 29190 21300 29294
rect 21420 29866 21540 31320
rect 22170 31110 22260 31320
rect 22410 31260 22950 31320
rect 22260 30990 22530 31110
rect 22740 31020 22860 31050
rect 21900 30495 22020 30510
rect 22140 30495 22260 30510
rect 21900 30480 22260 30495
rect 22440 30480 22530 30990
rect 21900 30405 22350 30480
rect 21900 30390 22020 30405
rect 22140 30390 22350 30405
rect 22440 30466 22590 30480
rect 22440 30390 22470 30466
rect 22260 30210 22350 30390
rect 21420 29280 21540 29294
rect 21660 29866 21780 29880
rect 21660 29190 21780 29294
rect 22230 29866 22350 29880
rect 22230 29190 22350 29294
rect 22470 29280 22590 29294
rect 22860 30466 22980 30480
rect 22860 29190 22980 29294
rect 23820 29880 23940 31605
rect 24780 31530 24990 31620
rect 25110 31906 25230 32010
rect 24060 31395 24180 31410
rect 24060 31305 24300 31395
rect 24060 31290 24180 31305
rect 24780 30210 24870 31530
rect 25110 31320 25230 31334
rect 25500 31906 25620 31920
rect 25980 31906 26100 31920
rect 25860 31605 25980 31695
rect 25500 31320 25620 31334
rect 25980 31320 26100 31334
rect 26220 31906 26340 31920
rect 26460 31890 26580 32010
rect 27420 31920 27540 32010
rect 26460 31440 26580 31470
rect 26700 31906 26820 31920
rect 26340 31334 26700 31350
rect 26220 31320 26820 31334
rect 25320 31230 25590 31320
rect 25320 31200 25410 31230
rect 25080 31110 25410 31200
rect 26010 31110 26100 31320
rect 26250 31260 26790 31320
rect 24780 30195 24900 30210
rect 24180 30105 24900 30195
rect 24780 30090 24900 30105
rect 24780 29880 24870 30090
rect 24990 30060 25080 31110
rect 25500 31095 25620 31110
rect 25500 31005 25740 31095
rect 25500 30990 25620 31005
rect 25980 30990 26370 31110
rect 26580 31020 26700 31050
rect 25170 30390 25260 30510
rect 25380 30405 25740 30495
rect 26280 30480 26370 30990
rect 26460 30795 26580 30810
rect 27180 30795 27300 31650
rect 27420 31620 27540 31650
rect 27750 31906 27870 31920
rect 27420 31290 27540 31410
rect 28140 31906 28260 32010
rect 27870 31334 28020 31410
rect 27750 31320 28020 31334
rect 28620 31920 28740 32010
rect 28620 31620 28740 31650
rect 28140 31320 28260 31334
rect 26460 30705 27300 30795
rect 26460 30690 26580 30705
rect 26100 30210 26190 30480
rect 26280 30466 26430 30480
rect 26280 30390 26310 30466
rect 24990 29970 25350 30060
rect 25260 29880 25350 29970
rect 23820 29280 23940 29310
rect 24060 29190 24180 29310
rect 24780 29866 24900 29880
rect 24780 29280 24900 29294
rect 25020 29866 25140 29880
rect 25020 29190 25140 29294
rect 25260 29866 25380 29880
rect 25260 29280 25380 29294
rect 25500 29866 25620 29880
rect 25500 29190 25620 29294
rect 26070 29866 26190 29880
rect 26070 29190 26190 29294
rect 26310 29280 26430 29294
rect 26700 30466 26820 30480
rect 26700 29190 26820 29294
rect 27180 29880 27300 30705
rect 27420 30495 27540 30510
rect 27660 30495 27780 30510
rect 27420 30405 27780 30495
rect 27420 30390 27540 30405
rect 27660 30390 27780 30405
rect 27180 29280 27300 29310
rect 27420 29190 27540 29310
rect 27660 29866 27780 29880
rect 27660 29190 27780 29294
rect 27900 29866 28020 31320
rect 28140 31095 28260 31110
rect 28140 31005 28380 31095
rect 28140 30990 28260 31005
rect 28860 30795 28980 31650
rect 29100 31906 29220 31920
rect 29100 31320 29220 31334
rect 29340 31906 29460 31920
rect 29580 31890 29700 32010
rect 29580 31440 29700 31470
rect 29820 31906 29940 31920
rect 29460 31334 29820 31350
rect 29340 31320 29940 31334
rect 30780 31906 30900 31920
rect 31020 31876 31170 32010
rect 31950 31920 32070 32010
rect 31020 31454 31034 31876
rect 31156 31454 31170 31876
rect 31020 31410 31170 31454
rect 31440 31860 31680 31920
rect 31440 31440 31500 31860
rect 31620 31440 31680 31860
rect 30780 31320 30900 31334
rect 31440 31380 31680 31440
rect 31950 31876 32100 31920
rect 31950 31454 31964 31876
rect 32086 31454 32100 31876
rect 31950 31410 32100 31454
rect 32220 31906 32340 31920
rect 29130 31110 29220 31320
rect 29370 31260 29910 31320
rect 30780 31230 31020 31320
rect 29100 30990 29490 31110
rect 31230 31110 31320 31170
rect 29700 31020 29820 31050
rect 30780 31095 30900 31110
rect 30180 31005 30900 31095
rect 30780 30990 30900 31005
rect 31440 31080 31530 31380
rect 32220 31320 32340 31334
rect 33180 31906 33300 32010
rect 33570 31906 33690 31920
rect 33180 31320 33300 31334
rect 32070 31230 32340 31320
rect 33540 31334 33570 31410
rect 33540 31320 33690 31334
rect 34620 31906 34740 32010
rect 35010 31906 35130 31920
rect 34620 31320 34740 31334
rect 34860 31334 35010 31410
rect 36060 31906 36180 31920
rect 35130 31334 35820 31395
rect 31440 30990 31590 31080
rect 32010 31050 32100 31080
rect 29100 30795 29220 30810
rect 28860 30705 29220 30795
rect 28860 29880 28980 30705
rect 29100 30690 29220 30705
rect 29400 30480 29490 30990
rect 29580 30690 29700 30810
rect 31500 30810 31590 30990
rect 31800 30960 32100 31050
rect 31500 30690 31620 30810
rect 31500 30480 31590 30690
rect 29220 30210 29310 30480
rect 29400 30466 29550 30480
rect 29400 30390 29430 30466
rect 27900 29280 28020 29294
rect 28140 29866 28260 29880
rect 28140 29190 28260 29294
rect 28620 29190 28740 29310
rect 28860 29280 28980 29310
rect 29190 29866 29310 29880
rect 29190 29190 29310 29294
rect 29430 29280 29550 29294
rect 29820 30466 29940 30480
rect 29820 29190 29940 29294
rect 30780 30466 31020 30480
rect 30900 30390 31020 30466
rect 31440 30466 31680 30480
rect 30780 29280 30900 29294
rect 31020 30210 31170 30270
rect 31020 29340 31034 30210
rect 31156 29340 31170 30210
rect 31020 29190 31170 29340
rect 31440 29294 31500 30466
rect 31620 29294 31680 30466
rect 32070 30466 32340 30480
rect 32070 30390 32220 30466
rect 31440 29280 31680 29294
rect 31950 30210 32100 30270
rect 31950 29340 31964 30210
rect 32086 29340 32100 30210
rect 31950 29280 32100 29340
rect 32220 29280 32340 29294
rect 33180 29866 33300 29880
rect 31950 29190 32070 29280
rect 33180 29190 33300 29294
rect 33420 29866 33540 31290
rect 34860 31305 35820 31334
rect 34620 31095 34740 31110
rect 34020 31005 34740 31095
rect 34620 30990 34740 31005
rect 33660 30390 33780 30510
rect 33420 29280 33540 29294
rect 33660 29866 33780 29880
rect 33660 29190 33780 29294
rect 34620 29866 34740 29880
rect 34620 29190 34740 29294
rect 34860 29866 34980 31305
rect 36060 31320 36180 31334
rect 36300 31906 36420 31920
rect 36540 31890 36660 32010
rect 36540 31440 36660 31470
rect 36780 31906 36900 31920
rect 36420 31334 36780 31350
rect 36300 31320 36900 31334
rect 37740 31906 37860 32010
rect 38130 31906 38250 31920
rect 37740 31320 37860 31334
rect 37980 31334 38130 31410
rect 37980 31320 38250 31334
rect 38940 31906 39060 31920
rect 39180 31890 39300 32010
rect 40860 31920 40980 32010
rect 39180 31440 39300 31470
rect 39420 31906 39540 31920
rect 39060 31334 39420 31350
rect 38940 31320 39540 31334
rect 39660 31906 39780 31920
rect 39660 31320 39780 31334
rect 36090 31110 36180 31320
rect 36330 31260 36870 31320
rect 36060 31095 36450 31110
rect 35220 31005 36450 31095
rect 36780 31050 36900 31110
rect 37740 31095 37860 31110
rect 36660 31020 36900 31050
rect 36060 30990 36450 31005
rect 36780 30990 36900 31020
rect 37035 31005 37860 31095
rect 35100 30390 35220 30510
rect 36060 30480 36180 30510
rect 36360 30480 36450 30990
rect 37035 30795 37125 31005
rect 37740 30990 37860 31005
rect 36660 30705 37125 30795
rect 36060 30390 36270 30480
rect 36360 30466 36510 30480
rect 36360 30390 36390 30466
rect 36180 30210 36270 30390
rect 34860 29280 34980 29294
rect 35100 29866 35220 29880
rect 35100 29190 35220 29294
rect 36150 29866 36270 29880
rect 36150 29190 36270 29294
rect 36390 29280 36510 29294
rect 36780 30466 36900 30480
rect 37980 30195 38100 31320
rect 38970 31260 39510 31320
rect 38940 31095 39060 31110
rect 38580 31050 39060 31095
rect 39660 31110 39750 31320
rect 38580 31020 39180 31050
rect 38580 31005 39060 31020
rect 38940 30990 39060 31005
rect 39390 30990 39780 31110
rect 39180 30690 39300 30810
rect 39390 30480 39480 30990
rect 39660 30795 39780 30810
rect 40620 30795 40740 31650
rect 40860 31620 40980 31650
rect 41670 31906 41790 31920
rect 40860 31395 40980 31410
rect 40860 31305 41340 31395
rect 40860 31290 40980 31305
rect 42060 31906 42180 32010
rect 41790 31334 41940 31410
rect 41670 31320 41940 31334
rect 42060 31320 42180 31334
rect 43020 31906 43140 31920
rect 43020 31320 43140 31334
rect 43260 31906 43380 31920
rect 43500 31890 43620 32010
rect 43500 31440 43620 31470
rect 43740 31906 43860 31920
rect 43380 31334 43740 31350
rect 43260 31320 43860 31334
rect 44460 31906 44580 31920
rect 44700 31890 44820 32010
rect 44700 31440 44820 31470
rect 44940 31906 45060 31920
rect 44580 31334 44940 31350
rect 44460 31320 45060 31334
rect 45180 31906 45300 31920
rect 46230 31906 46350 31920
rect 45300 31605 45660 31695
rect 45180 31320 45300 31334
rect 46620 31906 46740 32010
rect 48330 31920 48450 32010
rect 46350 31334 46500 31410
rect 46230 31320 46500 31334
rect 46620 31320 46740 31334
rect 48060 31906 48180 31920
rect 48300 31876 48450 31920
rect 48300 31454 48314 31876
rect 48436 31454 48450 31876
rect 48300 31410 48450 31454
rect 48720 31860 48960 31920
rect 48720 31440 48780 31860
rect 48900 31440 48960 31860
rect 48720 31380 48960 31440
rect 49230 31876 49380 32010
rect 49230 31454 49244 31876
rect 49366 31454 49380 31876
rect 49230 31410 49380 31454
rect 49500 31906 49620 31920
rect 48060 31320 48180 31334
rect 39660 30705 40740 30795
rect 39660 30690 39780 30705
rect 39660 30495 39780 30510
rect 40380 30495 40500 30510
rect 39660 30480 40500 30495
rect 38940 30466 39060 30480
rect 37620 30105 38100 30195
rect 36780 29190 36900 29294
rect 37740 29866 37860 29880
rect 37740 29190 37860 29294
rect 37980 29866 38100 30105
rect 37980 29280 38100 29294
rect 38220 29866 38340 29880
rect 38220 29190 38340 29294
rect 38940 29190 39060 29294
rect 39330 30466 39480 30480
rect 39450 30390 39480 30466
rect 39570 30405 40500 30480
rect 39570 30390 39780 30405
rect 40380 30390 40500 30405
rect 39570 30210 39660 30390
rect 40620 29880 40740 30705
rect 40980 30405 41580 30495
rect 41820 30495 41940 31320
rect 43050 31110 43140 31320
rect 43290 31260 43830 31320
rect 44490 31260 45030 31320
rect 42060 31095 42180 31110
rect 42780 31095 42900 31110
rect 42060 31005 42900 31095
rect 42060 30990 42180 31005
rect 42780 30990 42900 31005
rect 43020 30990 43260 31110
rect 43380 30990 43410 31110
rect 43620 31020 43740 31050
rect 44460 31095 44580 31110
rect 44100 31050 44580 31095
rect 45180 31110 45270 31320
rect 44100 31020 44700 31050
rect 44100 31005 44580 31020
rect 44460 30990 44580 31005
rect 44910 30990 45300 31110
rect 43020 30495 43140 30510
rect 41820 30480 43140 30495
rect 43320 30480 43410 30990
rect 44700 30795 44820 30810
rect 44100 30705 44820 30795
rect 44700 30690 44820 30705
rect 44910 30480 45000 30990
rect 46380 30795 46500 31320
rect 48060 31230 48330 31320
rect 48060 31095 48180 31110
rect 47460 31005 48180 31095
rect 48060 30990 48180 31005
rect 48870 31080 48960 31380
rect 49500 31320 49620 31334
rect 49380 31230 49620 31320
rect 48300 31050 48390 31080
rect 48300 30960 48600 31050
rect 48810 30990 48960 31080
rect 49080 31110 49170 31170
rect 49500 31095 49620 31110
rect 49500 31005 49740 31095
rect 49500 30990 49620 31005
rect 48810 30810 48900 30990
rect 45915 30705 46500 30795
rect 45180 30495 45300 30510
rect 45915 30495 46005 30705
rect 45180 30480 46005 30495
rect 41820 30405 43230 30480
rect 39330 29280 39450 29294
rect 39570 29866 39690 29880
rect 39570 29190 39690 29294
rect 40620 29280 40740 29310
rect 40860 29190 40980 29310
rect 41580 29866 41700 29880
rect 41580 29190 41700 29294
rect 41820 29866 41940 30405
rect 43020 30390 43230 30405
rect 43320 30466 43470 30480
rect 43320 30390 43350 30466
rect 43140 30210 43230 30390
rect 41820 29280 41940 29294
rect 42060 29866 42180 29880
rect 42060 29190 42180 29294
rect 43110 29866 43230 29880
rect 43110 29190 43230 29294
rect 43350 29280 43470 29294
rect 43740 30466 43860 30480
rect 43740 29190 43860 29294
rect 44460 30466 44580 30480
rect 44460 29190 44580 29294
rect 44850 30466 45000 30480
rect 44970 30390 45000 30466
rect 45090 30405 46005 30480
rect 45090 30390 45300 30405
rect 45090 30210 45180 30390
rect 44850 29280 44970 29294
rect 45090 29866 45210 29880
rect 45090 29190 45210 29294
rect 46140 29866 46260 29880
rect 46140 29190 46260 29294
rect 46380 29866 46500 30705
rect 48780 30795 48900 30810
rect 48780 30705 49500 30795
rect 48780 30690 48900 30705
rect 48810 30480 48900 30690
rect 48060 30466 48330 30480
rect 46380 29280 46500 29294
rect 46620 29866 46740 29880
rect 46620 29190 46740 29294
rect 48180 30390 48330 30466
rect 48720 30466 48960 30480
rect 48060 29280 48180 29294
rect 48300 30210 48450 30270
rect 48300 29340 48314 30210
rect 48436 29340 48450 30210
rect 48300 29280 48450 29340
rect 48720 29294 48780 30466
rect 48900 29294 48960 30466
rect 49380 30466 49620 30480
rect 49380 30390 49500 30466
rect 48720 29280 48960 29294
rect 49230 30210 49380 30270
rect 49230 29340 49244 30210
rect 49366 29340 49380 30210
rect 48330 29190 48450 29280
rect 49230 29190 49380 29340
rect 49500 29280 49620 29294
rect 1155 29160 54240 29190
rect 1155 29040 1214 29160
rect 2086 29040 5220 29160
rect 5340 29040 5460 29160
rect 5580 29040 5700 29160
rect 5820 29040 5940 29160
rect 6060 29040 6180 29160
rect 6300 29040 6420 29160
rect 6540 29040 6660 29160
rect 6780 29040 6900 29160
rect 7020 29040 7140 29160
rect 7260 29040 7380 29160
rect 7500 29040 7620 29160
rect 7740 29040 7860 29160
rect 7980 29040 8340 29160
rect 8460 29040 8580 29160
rect 8700 29040 8820 29160
rect 8940 29040 9060 29160
rect 9180 29040 9300 29160
rect 9420 29040 9540 29160
rect 9660 29040 9780 29160
rect 9900 29040 10020 29160
rect 10140 29040 10260 29160
rect 10380 29040 10500 29160
rect 10620 29040 10740 29160
rect 10860 29040 10980 29160
rect 11100 29040 11460 29160
rect 11580 29040 11940 29160
rect 12060 29040 12420 29160
rect 12540 29040 12660 29160
rect 12780 29040 12900 29160
rect 13020 29040 13140 29160
rect 13260 29040 13380 29160
rect 13500 29040 13620 29160
rect 13740 29040 13860 29160
rect 13980 29040 14100 29160
rect 14220 29040 14340 29160
rect 14460 29040 14580 29160
rect 14700 29040 14820 29160
rect 14940 29040 15060 29160
rect 15180 29040 15300 29160
rect 15420 29040 15540 29160
rect 15660 29040 15780 29160
rect 15900 29040 16020 29160
rect 16140 29040 16260 29160
rect 16380 29040 16500 29160
rect 16620 29040 16740 29160
rect 16860 29040 16980 29160
rect 17100 29040 17220 29160
rect 17340 29040 17460 29160
rect 17580 29040 17700 29160
rect 17820 29040 17940 29160
rect 18060 29040 18420 29160
rect 18540 29040 18660 29160
rect 18780 29040 18900 29160
rect 19020 29040 19140 29160
rect 19260 29040 19620 29160
rect 19740 29040 20100 29160
rect 20220 29040 20340 29160
rect 20460 29040 20580 29160
rect 20700 29040 20820 29160
rect 20940 29040 21060 29160
rect 21180 29040 21300 29160
rect 21420 29040 21540 29160
rect 21660 29040 21780 29160
rect 21900 29040 22020 29160
rect 22140 29040 22500 29160
rect 22620 29040 22740 29160
rect 22860 29040 22980 29160
rect 23100 29040 23220 29160
rect 23340 29040 23460 29160
rect 23580 29040 23700 29160
rect 23820 29040 23940 29160
rect 24060 29040 24180 29160
rect 24300 29040 24420 29160
rect 24540 29040 24660 29160
rect 24780 29040 24900 29160
rect 25020 29040 25140 29160
rect 25260 29040 25380 29160
rect 25500 29040 25620 29160
rect 25740 29040 25860 29160
rect 25980 29040 26100 29160
rect 26220 29040 26340 29160
rect 26460 29040 26820 29160
rect 26940 29040 27060 29160
rect 27180 29040 27300 29160
rect 27420 29040 27540 29160
rect 27660 29040 27780 29160
rect 27900 29040 28020 29160
rect 28140 29040 28260 29160
rect 28380 29040 28500 29160
rect 28620 29040 28740 29160
rect 28860 29040 29220 29160
rect 29340 29040 29460 29160
rect 29580 29040 29700 29160
rect 29820 29040 29940 29160
rect 30060 29040 30180 29160
rect 30300 29040 30420 29160
rect 30540 29040 30660 29160
rect 30780 29040 30900 29160
rect 31020 29040 31140 29160
rect 31260 29040 31380 29160
rect 31500 29040 31620 29160
rect 31740 29040 31860 29160
rect 31980 29040 32100 29160
rect 32220 29040 32340 29160
rect 32460 29040 32580 29160
rect 32700 29040 32820 29160
rect 32940 29040 33060 29160
rect 33180 29040 33300 29160
rect 33420 29040 33540 29160
rect 33660 29040 33780 29160
rect 33900 29040 34020 29160
rect 34140 29040 34260 29160
rect 34380 29040 34500 29160
rect 34620 29040 34740 29160
rect 34860 29040 34980 29160
rect 35100 29040 35220 29160
rect 35340 29040 35460 29160
rect 35580 29040 35700 29160
rect 35820 29040 35940 29160
rect 36060 29040 36420 29160
rect 36540 29040 36660 29160
rect 36780 29040 36900 29160
rect 37020 29040 37140 29160
rect 37260 29040 37380 29160
rect 37500 29040 37620 29160
rect 37740 29040 38100 29160
rect 38220 29040 38340 29160
rect 38460 29040 38580 29160
rect 38700 29040 38820 29160
rect 38940 29040 39060 29160
rect 39180 29040 39300 29160
rect 39420 29040 39540 29160
rect 39660 29040 39780 29160
rect 39900 29040 40020 29160
rect 40140 29040 40260 29160
rect 40380 29040 40500 29160
rect 40620 29040 40980 29160
rect 41100 29040 41220 29160
rect 41340 29040 41460 29160
rect 41580 29040 41700 29160
rect 41820 29040 41940 29160
rect 42060 29040 42180 29160
rect 42300 29040 42420 29160
rect 42540 29040 42660 29160
rect 42780 29040 42900 29160
rect 43020 29040 43380 29160
rect 43500 29040 43860 29160
rect 43980 29040 44100 29160
rect 44220 29040 44340 29160
rect 44460 29040 44820 29160
rect 44940 29040 45300 29160
rect 45420 29040 45540 29160
rect 45660 29040 45780 29160
rect 45900 29040 46020 29160
rect 46140 29040 46260 29160
rect 46380 29040 46740 29160
rect 46860 29040 46980 29160
rect 47100 29040 47220 29160
rect 47340 29040 47460 29160
rect 47580 29040 47700 29160
rect 47820 29040 47940 29160
rect 48060 29040 48420 29160
rect 48540 29040 48900 29160
rect 49020 29040 49140 29160
rect 49260 29040 49380 29160
rect 49500 29040 49620 29160
rect 49740 29040 49860 29160
rect 49980 29040 50100 29160
rect 50220 29040 53310 29160
rect 54180 29040 54240 29160
rect 1155 29010 54240 29040
rect 7290 28920 7410 29010
rect 7020 28906 7140 28920
rect 7260 28860 7410 28920
rect 7260 27990 7274 28860
rect 7396 27990 7410 28860
rect 7260 27930 7410 27990
rect 7680 28906 7920 28920
rect 7140 27734 7290 27810
rect 7020 27720 7290 27734
rect 7680 27734 7740 28906
rect 7860 27734 7920 28906
rect 8190 28860 8340 29010
rect 8190 27990 8204 28860
rect 8326 27990 8340 28860
rect 8190 27930 8340 27990
rect 8460 28906 8580 28920
rect 7680 27720 7920 27734
rect 8340 27734 8460 27810
rect 8700 28906 8820 29010
rect 8700 28320 8820 28334
rect 8940 28906 9060 28920
rect 8340 27720 8580 27734
rect 7770 27510 7860 27720
rect 7740 27495 7860 27510
rect 8700 27495 8820 27510
rect 7740 27405 8820 27495
rect 7740 27390 7860 27405
rect 8700 27390 8820 27405
rect 7260 27150 7560 27240
rect 7770 27210 7860 27390
rect 7260 27120 7350 27150
rect 7770 27120 7920 27210
rect 7020 26880 7290 26970
rect 7020 26866 7140 26880
rect 7830 26820 7920 27120
rect 8040 27030 8130 27090
rect 8340 26880 8580 26970
rect 8940 26880 9060 28334
rect 9180 28906 9300 29010
rect 9180 28320 9300 28334
rect 9420 28906 9540 28920
rect 9660 28860 9810 29010
rect 10590 28920 10710 29010
rect 9660 27990 9674 28860
rect 9796 27990 9810 28860
rect 9660 27930 9810 27990
rect 10080 28906 10320 28920
rect 9540 27734 9660 27810
rect 9420 27720 9660 27734
rect 10080 27810 10140 28906
rect 10020 27734 10140 27810
rect 10260 27734 10320 28906
rect 10590 28860 10740 28920
rect 10590 27990 10604 28860
rect 10726 27990 10740 28860
rect 10590 27930 10740 27990
rect 10860 28906 10980 28920
rect 10020 27720 10320 27734
rect 10770 27734 10860 27810
rect 10770 27720 10980 27734
rect 11100 28906 11220 29010
rect 11100 27720 11220 27734
rect 11490 28906 11610 28920
rect 11730 28906 11850 29010
rect 11730 28320 11850 28334
rect 12060 28906 12180 29010
rect 12060 28320 12180 28334
rect 12300 28906 12420 28920
rect 11730 27810 11820 27990
rect 11610 27734 11640 27810
rect 11490 27720 11640 27734
rect 11730 27795 11940 27810
rect 12300 27795 12420 28334
rect 12540 28906 12660 29010
rect 12540 28320 12660 28334
rect 12780 28906 12900 29010
rect 12780 28320 12900 28334
rect 13020 28906 13140 28920
rect 11730 27720 12420 27795
rect 10020 27510 10110 27720
rect 10650 27630 10740 27720
rect 10350 27540 10740 27630
rect 9900 27420 10110 27510
rect 9900 27390 10170 27420
rect 10020 27330 10170 27390
rect 9420 27195 9540 27210
rect 9300 27105 9540 27195
rect 9420 27090 9540 27105
rect 9870 27030 9960 27090
rect 9420 26880 9660 26970
rect 7020 26280 7140 26294
rect 7260 26746 7410 26790
rect 7260 26324 7274 26746
rect 7396 26324 7410 26746
rect 7260 26280 7410 26324
rect 7680 26760 7920 26820
rect 8460 26866 8580 26880
rect 7680 26340 7740 26760
rect 7860 26340 7920 26760
rect 7680 26280 7920 26340
rect 8190 26746 8340 26790
rect 8190 26324 8204 26746
rect 8326 26324 8340 26746
rect 7290 26190 7410 26280
rect 8190 26190 8340 26324
rect 8460 26280 8580 26294
rect 8700 26866 8820 26880
rect 8940 26866 9210 26880
rect 8940 26790 9090 26866
rect 8700 26190 8820 26294
rect 9090 26280 9210 26294
rect 9420 26866 9540 26880
rect 10080 26820 10170 27330
rect 10290 27330 10560 27420
rect 10290 27240 10380 27330
rect 11550 27210 11640 27720
rect 11820 27705 12420 27720
rect 11820 27690 11940 27705
rect 10470 27090 10740 27180
rect 10860 27090 10980 27210
rect 11100 27180 11220 27210
rect 11100 27150 11340 27180
rect 11100 27090 11220 27150
rect 10470 27030 10560 27090
rect 11550 27090 11820 27210
rect 10500 26940 10560 27030
rect 10770 26880 10980 26970
rect 11130 26880 11670 26940
rect 11820 26880 11910 27090
rect 12300 26880 12420 27705
rect 12540 27795 12660 27810
rect 13020 27795 13140 28334
rect 13260 28906 13380 29010
rect 13260 28320 13380 28334
rect 13740 28906 13860 28920
rect 13740 28320 13860 28334
rect 13980 28906 14100 29010
rect 13980 28320 14100 28334
rect 14220 28906 14340 28920
rect 14220 28320 14340 28334
rect 14460 28906 14580 29010
rect 14460 28320 14580 28334
rect 15420 28906 15540 29010
rect 15420 28320 15540 28334
rect 15660 28906 15780 28920
rect 13740 28110 13830 28320
rect 14220 28230 14310 28320
rect 13950 28140 14310 28230
rect 13740 27990 13860 28110
rect 12540 27705 13140 27795
rect 12540 27690 12660 27705
rect 12540 27195 12660 27210
rect 12780 27195 12900 27210
rect 12540 27105 12900 27195
rect 12540 27090 12660 27105
rect 12780 27090 12900 27105
rect 13020 26880 13140 27705
rect 13260 27690 13380 27810
rect 10860 26866 10980 26880
rect 9420 26280 9540 26294
rect 9660 26746 9810 26790
rect 9660 26324 9674 26746
rect 9796 26324 9810 26746
rect 9660 26190 9810 26324
rect 10080 26760 10320 26820
rect 10080 26340 10140 26760
rect 10260 26340 10320 26760
rect 10080 26280 10320 26340
rect 10590 26746 10740 26790
rect 10590 26324 10604 26746
rect 10726 26324 10740 26746
rect 10590 26280 10740 26324
rect 10860 26280 10980 26294
rect 11100 26866 11700 26880
rect 11220 26850 11580 26866
rect 11100 26280 11220 26294
rect 11340 26730 11460 26760
rect 10590 26190 10710 26280
rect 11340 26190 11460 26310
rect 11580 26280 11700 26294
rect 11820 26866 11940 26880
rect 11820 26280 11940 26294
rect 12060 26866 12180 26880
rect 12300 26866 12570 26880
rect 12300 26790 12450 26866
rect 12060 26190 12180 26294
rect 12450 26280 12570 26294
rect 12780 26866 12900 26880
rect 13020 26866 13290 26880
rect 13020 26790 13170 26866
rect 12780 26190 12900 26294
rect 13740 26670 13830 27990
rect 13950 27090 14040 28140
rect 15660 28095 15780 28334
rect 15900 28906 16020 29010
rect 15900 28320 16020 28334
rect 16620 28906 16740 29010
rect 16620 28320 16740 28334
rect 16860 28906 16980 28920
rect 14580 28005 15780 28095
rect 14130 27795 14340 27810
rect 15180 27795 15300 27810
rect 14130 27705 15300 27795
rect 14130 27690 14340 27705
rect 15180 27690 15300 27705
rect 14460 27195 14580 27210
rect 14460 27105 15180 27195
rect 14460 27090 14580 27105
rect 14040 27000 14370 27090
rect 14280 26970 14370 27000
rect 14280 26880 14550 26970
rect 15660 26880 15780 28005
rect 15900 27795 16020 27810
rect 15900 27705 16380 27795
rect 15900 27690 16020 27705
rect 16500 27705 16620 27795
rect 16860 26880 16980 28334
rect 17100 28906 17220 29010
rect 17100 28320 17220 28334
rect 18060 28906 18180 29010
rect 18060 28320 18180 28334
rect 18300 28906 18420 28920
rect 17100 27195 17220 27210
rect 17100 27105 17820 27195
rect 17100 27090 17220 27105
rect 18060 27090 18180 27210
rect 18300 26910 18420 28334
rect 18540 28906 18660 29010
rect 18540 28320 18660 28334
rect 19350 28906 19470 29010
rect 19350 28320 19470 28334
rect 19590 28906 19710 28920
rect 18540 27795 18660 27810
rect 18540 27705 18780 27795
rect 18540 27690 18660 27705
rect 19380 27720 19470 27990
rect 19560 27734 19590 27810
rect 19560 27720 19710 27734
rect 19980 28906 20100 29010
rect 20940 28906 21060 29010
rect 20940 28320 21060 28334
rect 21180 28906 21300 28920
rect 19980 27720 20100 27734
rect 19560 27210 19650 27720
rect 19260 27090 19650 27210
rect 19980 27195 20100 27210
rect 20700 27195 20820 27210
rect 19980 27180 20820 27195
rect 19860 27150 20820 27180
rect 14070 26866 14190 26880
rect 13740 26580 13950 26670
rect 13170 26280 13290 26294
rect 13830 26566 13950 26580
rect 13830 26280 13950 26294
rect 14070 26190 14190 26294
rect 14460 26866 14580 26880
rect 14460 26280 14580 26294
rect 15420 26866 15540 26880
rect 15660 26866 15930 26880
rect 15660 26790 15810 26866
rect 15420 26190 15540 26294
rect 15810 26280 15930 26294
rect 16710 26866 16980 26880
rect 16830 26790 16980 26866
rect 17100 26866 17220 26880
rect 16710 26280 16830 26294
rect 17100 26190 17220 26294
rect 18060 26866 18180 26880
rect 19290 26880 19380 27090
rect 19980 27105 20820 27150
rect 19980 27090 20100 27105
rect 20700 27090 20820 27105
rect 19530 26880 20070 26940
rect 21180 26880 21300 28334
rect 21420 28906 21540 29010
rect 21420 28320 21540 28334
rect 22140 28906 22260 29010
rect 22140 28320 22260 28334
rect 22380 28906 22500 28920
rect 21660 28095 21780 28110
rect 22380 28095 22500 28334
rect 22620 28906 22740 29010
rect 22620 28320 22740 28334
rect 23580 28906 23700 29010
rect 23580 28320 23700 28334
rect 23820 28906 23940 28920
rect 21660 28005 22500 28095
rect 21660 27990 21780 28005
rect 22140 27195 22260 27210
rect 21780 27105 22260 27195
rect 22140 27090 22260 27105
rect 22380 26880 22500 28005
rect 23820 28095 23940 28334
rect 24060 28906 24180 29010
rect 24060 28320 24180 28334
rect 25020 28906 25140 29010
rect 25020 28320 25140 28334
rect 25260 28906 25380 28920
rect 22980 28005 23940 28095
rect 22620 27795 22740 27810
rect 22620 27705 23580 27795
rect 22620 27690 22740 27705
rect 23220 27105 23580 27195
rect 23820 26880 23940 28005
rect 24060 27690 24180 27810
rect 25020 27195 25140 27210
rect 24180 27105 25140 27195
rect 25020 27090 25140 27105
rect 25260 26880 25380 28334
rect 25500 28906 25620 29010
rect 25500 28320 25620 28334
rect 26460 28906 26580 29010
rect 26460 28320 26580 28334
rect 26700 28906 26820 28920
rect 26700 27495 26820 28334
rect 26940 28906 27060 29010
rect 26940 28320 27060 28334
rect 28470 28906 28590 29010
rect 28470 28320 28590 28334
rect 28710 28906 28830 28920
rect 28500 27810 28590 27990
rect 26940 27795 27060 27810
rect 26940 27705 27180 27795
rect 26940 27690 27060 27705
rect 28380 27795 28590 27810
rect 28020 27720 28590 27795
rect 28680 27734 28710 27810
rect 28680 27720 28830 27734
rect 29100 28906 29220 29010
rect 30300 28906 30420 29010
rect 30300 28320 30420 28334
rect 30540 28906 30660 28920
rect 29100 27720 29220 27734
rect 28020 27705 28500 27720
rect 28380 27690 28500 27705
rect 28380 27495 28500 27510
rect 26700 27405 28500 27495
rect 26460 27195 26580 27210
rect 25620 27105 26580 27195
rect 26460 27090 26580 27105
rect 26700 26880 26820 27405
rect 28380 27390 28500 27405
rect 28680 27210 28770 27720
rect 29460 27705 30300 27795
rect 30540 27795 30660 28334
rect 30780 28906 30900 29010
rect 30780 28320 30900 28334
rect 31830 28906 31950 29010
rect 31830 28320 31950 28334
rect 32070 28906 32190 28920
rect 31860 27810 31950 27990
rect 31740 27795 31950 27810
rect 30540 27720 31950 27795
rect 32040 27734 32070 27810
rect 32040 27720 32190 27734
rect 32460 28906 32580 29010
rect 33210 28920 33330 29010
rect 32460 27720 32580 27734
rect 32940 28906 33060 28920
rect 33180 28860 33330 28920
rect 33180 27990 33194 28860
rect 33316 27990 33330 28860
rect 33180 27930 33330 27990
rect 33600 28906 33840 28920
rect 33060 27734 33210 27810
rect 32940 27720 33210 27734
rect 33600 27734 33660 28906
rect 33780 27734 33840 28906
rect 34110 28860 34260 29010
rect 34110 27990 34124 28860
rect 34246 27990 34260 28860
rect 34110 27930 34260 27990
rect 34380 28906 34500 28920
rect 33600 27720 33840 27734
rect 34260 27734 34380 27810
rect 34860 28906 34980 29010
rect 34860 28320 34980 28334
rect 35100 28906 35220 28920
rect 34260 27720 34500 27734
rect 30540 27705 31860 27720
rect 28860 27390 28980 27510
rect 28380 27090 28620 27210
rect 28740 27090 28770 27210
rect 28980 27150 29100 27180
rect 28410 26880 28500 27090
rect 28650 26880 29190 26940
rect 30540 26880 30660 27705
rect 31740 27690 31860 27705
rect 32040 27210 32130 27720
rect 32220 27390 32340 27510
rect 33690 27510 33780 27720
rect 33660 27390 33780 27510
rect 31740 27090 32130 27210
rect 32340 27150 32460 27180
rect 31770 26880 31860 27090
rect 32940 27195 33060 27210
rect 32820 27105 33060 27195
rect 32940 27090 33060 27105
rect 33180 27150 33480 27240
rect 33690 27210 33780 27390
rect 33180 27120 33270 27150
rect 33690 27120 33840 27210
rect 32010 26880 32550 26940
rect 32940 26880 33210 26970
rect 18420 26866 18570 26880
rect 18420 26790 18450 26866
rect 18060 26190 18180 26294
rect 19260 26866 19380 26880
rect 18900 26505 19260 26595
rect 18450 26280 18570 26294
rect 19260 26280 19380 26294
rect 19500 26866 20100 26880
rect 19620 26850 19980 26866
rect 19500 26280 19620 26294
rect 19740 26730 19860 26760
rect 19740 26190 19860 26310
rect 19980 26280 20100 26294
rect 20940 26866 21060 26880
rect 21180 26866 21450 26880
rect 21180 26790 21330 26866
rect 20940 26190 21060 26294
rect 21330 26280 21450 26294
rect 22140 26866 22260 26880
rect 22380 26866 22650 26880
rect 22380 26790 22530 26866
rect 22140 26190 22260 26294
rect 22530 26280 22650 26294
rect 23580 26866 23700 26880
rect 23820 26866 24090 26880
rect 23820 26790 23970 26866
rect 23580 26190 23700 26294
rect 23970 26280 24090 26294
rect 25020 26866 25140 26880
rect 25260 26866 25530 26880
rect 25260 26790 25410 26866
rect 25020 26190 25140 26294
rect 25410 26280 25530 26294
rect 26460 26866 26580 26880
rect 26700 26866 26970 26880
rect 26700 26790 26850 26866
rect 26460 26190 26580 26294
rect 26850 26280 26970 26294
rect 28380 26866 28500 26880
rect 28380 26280 28500 26294
rect 28620 26866 29220 26880
rect 28740 26850 29100 26866
rect 28620 26280 28740 26294
rect 28860 26730 28980 26760
rect 28860 26190 28980 26310
rect 29100 26280 29220 26294
rect 30390 26866 30660 26880
rect 30510 26790 30660 26866
rect 30780 26866 30900 26880
rect 30390 26280 30510 26294
rect 30780 26190 30900 26294
rect 31740 26866 31860 26880
rect 31740 26280 31860 26294
rect 31980 26866 32580 26880
rect 32100 26850 32460 26866
rect 31980 26280 32100 26294
rect 32220 26730 32340 26760
rect 32220 26190 32340 26310
rect 32460 26280 32580 26294
rect 32940 26866 33060 26880
rect 33750 26820 33840 27120
rect 34380 27090 34500 27210
rect 34860 27195 34980 27210
rect 34740 27105 34980 27195
rect 34860 27090 34980 27105
rect 33960 27030 34050 27090
rect 34260 26880 34500 26970
rect 35100 26880 35220 28334
rect 35340 28906 35460 29010
rect 35340 28320 35460 28334
rect 36060 28906 36180 29010
rect 36060 28320 36180 28334
rect 36300 28906 36420 28920
rect 36060 27195 36180 27210
rect 35700 27105 36180 27195
rect 36060 27090 36180 27105
rect 36300 26880 36420 28334
rect 36540 28906 36660 29010
rect 36540 28320 36660 28334
rect 37500 28906 37620 29010
rect 37500 28320 37620 28334
rect 37740 28906 37860 28920
rect 36540 27795 36660 27810
rect 36540 27705 37020 27795
rect 36540 27690 36660 27705
rect 37140 27705 37260 27795
rect 37740 26880 37860 28334
rect 37980 28906 38100 29010
rect 37980 28320 38100 28334
rect 38700 28906 38820 29010
rect 38700 28320 38820 28334
rect 38940 28906 39060 28920
rect 37980 27195 38100 27210
rect 38460 27195 38580 27210
rect 37980 27105 38580 27195
rect 37980 27090 38100 27105
rect 38460 27090 38580 27105
rect 38940 26880 39060 28334
rect 39180 28906 39300 29010
rect 39930 28920 40050 29010
rect 39180 28320 39300 28334
rect 39660 28906 39780 28920
rect 39180 27795 39300 27810
rect 39180 27705 39420 27795
rect 39180 27690 39300 27705
rect 39900 28860 40050 28920
rect 39900 27990 39914 28860
rect 40036 27990 40050 28860
rect 39900 27930 40050 27990
rect 40320 28906 40560 28920
rect 39780 27734 39930 27810
rect 39660 27720 39930 27734
rect 40320 27734 40380 28906
rect 40500 27734 40560 28906
rect 40830 28860 40980 29010
rect 40830 27990 40844 28860
rect 40966 27990 40980 28860
rect 40830 27930 40980 27990
rect 41100 28906 41220 28920
rect 40320 27720 40560 27734
rect 40980 27734 41100 27810
rect 41580 28906 41700 29010
rect 41580 28320 41700 28334
rect 41820 28906 41940 28920
rect 40980 27720 41220 27734
rect 40410 27510 40500 27720
rect 40380 27390 40500 27510
rect 39660 27195 39780 27210
rect 39300 27105 39780 27195
rect 39660 27090 39780 27105
rect 39900 27150 40200 27240
rect 40410 27210 40500 27390
rect 41820 27495 41940 28334
rect 42060 28906 42180 29010
rect 42060 28320 42180 28334
rect 43110 28906 43230 29010
rect 43110 28320 43230 28334
rect 43350 28906 43470 28920
rect 43140 27810 43230 27990
rect 43020 27795 43230 27810
rect 42315 27720 43230 27795
rect 43320 27734 43350 27810
rect 43320 27720 43470 27734
rect 43740 28906 43860 29010
rect 43740 27720 43860 27734
rect 44460 28906 44580 29010
rect 44460 27720 44580 27734
rect 44850 28906 44970 28920
rect 45090 28906 45210 29010
rect 45090 28320 45210 28334
rect 45900 28906 46020 29010
rect 44970 27734 45000 27810
rect 44850 27720 45000 27734
rect 45090 27720 45180 27990
rect 42315 27705 43140 27720
rect 42315 27495 42405 27705
rect 43020 27690 43140 27705
rect 41820 27405 42405 27495
rect 39900 27120 39990 27150
rect 40410 27120 40560 27210
rect 39660 26880 39930 26970
rect 32940 26280 33060 26294
rect 33180 26746 33330 26790
rect 33180 26324 33194 26746
rect 33316 26324 33330 26746
rect 33180 26280 33330 26324
rect 33600 26760 33840 26820
rect 34380 26866 34500 26880
rect 33600 26340 33660 26760
rect 33780 26340 33840 26760
rect 33600 26280 33840 26340
rect 34110 26746 34260 26790
rect 34110 26324 34124 26746
rect 34246 26324 34260 26746
rect 33210 26190 33330 26280
rect 34110 26190 34260 26324
rect 34380 26280 34500 26294
rect 34860 26866 34980 26880
rect 35100 26866 35370 26880
rect 35100 26790 35250 26866
rect 34860 26190 34980 26294
rect 35250 26280 35370 26294
rect 36060 26866 36180 26880
rect 36300 26866 36570 26880
rect 36300 26790 36450 26866
rect 36060 26190 36180 26294
rect 36450 26280 36570 26294
rect 37590 26866 37860 26880
rect 37710 26790 37860 26866
rect 37980 26866 38100 26880
rect 37590 26280 37710 26294
rect 37980 26190 38100 26294
rect 38700 26866 38820 26880
rect 38940 26866 39210 26880
rect 38940 26790 39090 26866
rect 38700 26190 38820 26294
rect 39090 26280 39210 26294
rect 39660 26866 39780 26880
rect 40470 26820 40560 27120
rect 41340 27195 41460 27210
rect 41580 27195 41700 27210
rect 41340 27105 41700 27195
rect 41340 27090 41460 27105
rect 41580 27090 41700 27105
rect 40680 27030 40770 27090
rect 40980 26880 41220 26970
rect 41820 26880 41940 27405
rect 43320 27210 43410 27720
rect 44910 27210 45000 27720
rect 45900 27720 46020 27734
rect 46290 28906 46410 28920
rect 46530 28906 46650 29010
rect 46530 28320 46650 28334
rect 46860 28890 46980 29010
rect 48060 28920 48180 29010
rect 47100 28890 47220 28920
rect 46530 27810 46620 27990
rect 46410 27734 46440 27810
rect 46290 27720 46440 27734
rect 46530 27720 46740 27810
rect 46350 27210 46440 27720
rect 46620 27690 46740 27720
rect 43020 27195 43410 27210
rect 42900 27105 43410 27195
rect 43020 27090 43410 27105
rect 43620 27150 43740 27180
rect 43050 26880 43140 27090
rect 44580 27150 44700 27180
rect 44910 27090 44940 27210
rect 45060 27090 45300 27210
rect 46350 27195 46740 27210
rect 46860 27195 46980 27210
rect 46020 27150 46140 27180
rect 43290 26880 43830 26940
rect 44490 26880 45030 26940
rect 45180 26880 45270 27090
rect 46350 27105 46980 27195
rect 46350 27090 46740 27105
rect 46860 27090 46980 27105
rect 47100 27195 47220 28320
rect 47340 28906 47940 28920
rect 47460 28830 47820 28906
rect 47340 27720 47460 27734
rect 48300 28876 48420 28920
rect 48540 28906 48660 29010
rect 48540 28320 48660 28334
rect 48780 28906 48900 28920
rect 48300 27810 48420 27854
rect 47940 27734 48420 27810
rect 47820 27720 48420 27734
rect 47610 27630 47700 27720
rect 47610 27540 47910 27630
rect 47820 27510 47910 27540
rect 47820 27390 47940 27510
rect 48300 27450 48420 27510
rect 48180 27420 48420 27450
rect 48300 27390 48420 27420
rect 47610 27210 47700 27270
rect 47580 27195 47700 27210
rect 47100 27105 47700 27195
rect 45930 26880 46470 26940
rect 46620 26880 46710 27090
rect 39660 26280 39780 26294
rect 39900 26746 40050 26790
rect 39900 26324 39914 26746
rect 40036 26324 40050 26746
rect 39900 26280 40050 26324
rect 40320 26760 40560 26820
rect 41100 26866 41220 26880
rect 40320 26340 40380 26760
rect 40500 26340 40560 26760
rect 40320 26280 40560 26340
rect 40830 26746 40980 26790
rect 40830 26324 40844 26746
rect 40966 26324 40980 26746
rect 39930 26190 40050 26280
rect 40830 26190 40980 26324
rect 41100 26280 41220 26294
rect 41580 26866 41700 26880
rect 41820 26866 42090 26880
rect 41820 26790 41970 26866
rect 41580 26190 41700 26294
rect 41970 26280 42090 26294
rect 43020 26866 43140 26880
rect 43020 26280 43140 26294
rect 43260 26866 43860 26880
rect 43380 26850 43740 26866
rect 43260 26280 43380 26294
rect 43500 26730 43620 26760
rect 43500 26190 43620 26310
rect 43740 26280 43860 26294
rect 44460 26866 45060 26880
rect 44580 26850 44940 26866
rect 44460 26280 44580 26294
rect 44700 26730 44820 26760
rect 44700 26190 44820 26310
rect 44940 26280 45060 26294
rect 45180 26866 45300 26880
rect 45180 26280 45300 26294
rect 45900 26866 46500 26880
rect 46020 26850 46380 26866
rect 45900 26280 46020 26294
rect 46140 26730 46260 26760
rect 46140 26190 46260 26310
rect 46380 26280 46500 26294
rect 46620 26866 46740 26880
rect 46860 26790 46980 26910
rect 46620 26280 46740 26294
rect 46860 26550 46980 26580
rect 47100 26550 47220 27105
rect 47580 27090 47700 27105
rect 47820 26880 47910 27390
rect 48060 27090 48180 27210
rect 48315 27195 48405 27390
rect 48315 27105 48540 27195
rect 48780 26880 48900 28334
rect 49020 28906 49140 29010
rect 49020 28320 49140 28334
rect 49260 28906 49380 29010
rect 49260 27720 49380 27734
rect 49650 28906 49770 28920
rect 49890 28906 50010 29010
rect 49890 28320 50010 28334
rect 49890 27810 49980 27990
rect 49770 27734 49800 27810
rect 49650 27720 49800 27734
rect 49890 27720 50100 27810
rect 49020 27495 49140 27510
rect 49500 27495 49620 27510
rect 49020 27405 49620 27495
rect 49020 27390 49140 27405
rect 49500 27390 49620 27405
rect 49710 27210 49800 27720
rect 49980 27690 50100 27720
rect 49140 27105 49260 27195
rect 49380 27150 49500 27180
rect 49710 27090 49740 27210
rect 49860 27090 50100 27210
rect 49290 26880 49830 26940
rect 49980 26880 50070 27090
rect 47340 26866 47460 26880
rect 46860 26190 46980 26280
rect 47340 26190 47460 26294
rect 47730 26866 47970 26880
rect 47730 26294 47790 26866
rect 47910 26294 47970 26866
rect 47730 26280 47970 26294
rect 48240 26866 48360 26880
rect 48240 26190 48360 26294
rect 48540 26866 48660 26880
rect 48780 26866 49050 26880
rect 48780 26790 48930 26866
rect 48540 26190 48660 26294
rect 48930 26280 49050 26294
rect 49260 26866 49860 26880
rect 49380 26850 49740 26866
rect 49260 26280 49380 26294
rect 49500 26730 49620 26760
rect 49500 26190 49620 26310
rect 49740 26280 49860 26294
rect 49980 26866 50100 26880
rect 49980 26280 50100 26294
rect 3135 26160 52260 26190
rect 3135 26040 3194 26160
rect 4066 26040 5220 26160
rect 5340 26040 5460 26160
rect 5580 26040 5700 26160
rect 5820 26040 5940 26160
rect 6060 26040 6180 26160
rect 6300 26040 6420 26160
rect 6540 26040 6660 26160
rect 6780 26040 6900 26160
rect 7020 26040 7380 26160
rect 7500 26040 7860 26160
rect 7980 26040 8100 26160
rect 8220 26040 8340 26160
rect 8460 26040 8580 26160
rect 8700 26040 9060 26160
rect 9180 26040 9300 26160
rect 9420 26040 9540 26160
rect 9660 26040 9780 26160
rect 9900 26040 10020 26160
rect 10140 26040 10260 26160
rect 10380 26040 10500 26160
rect 10620 26040 10740 26160
rect 10860 26040 10980 26160
rect 11100 26040 11220 26160
rect 11340 26040 11460 26160
rect 11580 26040 11700 26160
rect 11820 26040 11940 26160
rect 12060 26040 12420 26160
rect 12540 26040 12660 26160
rect 12780 26040 12900 26160
rect 13020 26040 13140 26160
rect 13260 26040 13380 26160
rect 13500 26040 13620 26160
rect 13740 26040 14100 26160
rect 14220 26040 14340 26160
rect 14460 26040 14580 26160
rect 14700 26040 14820 26160
rect 14940 26040 15060 26160
rect 15180 26040 15300 26160
rect 15420 26040 15780 26160
rect 15900 26040 16020 26160
rect 16140 26040 16260 26160
rect 16380 26040 16500 26160
rect 16620 26040 16740 26160
rect 16860 26040 16980 26160
rect 17100 26040 17220 26160
rect 17340 26040 17460 26160
rect 17580 26040 17700 26160
rect 17820 26040 17940 26160
rect 18060 26040 18180 26160
rect 18300 26040 18420 26160
rect 18540 26040 18660 26160
rect 18780 26040 18900 26160
rect 19020 26040 19140 26160
rect 19260 26040 19380 26160
rect 19500 26040 19620 26160
rect 19740 26040 19860 26160
rect 19980 26040 20100 26160
rect 20220 26040 20340 26160
rect 20460 26040 20580 26160
rect 20700 26040 20820 26160
rect 20940 26040 21300 26160
rect 21420 26040 21540 26160
rect 21660 26040 21780 26160
rect 21900 26040 22020 26160
rect 22140 26040 22260 26160
rect 22380 26040 22500 26160
rect 22620 26040 22740 26160
rect 22860 26040 22980 26160
rect 23100 26040 23220 26160
rect 23340 26040 23460 26160
rect 23580 26040 23700 26160
rect 23820 26040 23940 26160
rect 24060 26040 24180 26160
rect 24300 26040 24420 26160
rect 24540 26040 24660 26160
rect 24780 26040 24900 26160
rect 25020 26040 25140 26160
rect 25260 26040 25380 26160
rect 25500 26040 25620 26160
rect 25740 26040 25860 26160
rect 25980 26040 26100 26160
rect 26220 26040 26340 26160
rect 26460 26040 26580 26160
rect 26700 26040 26820 26160
rect 26940 26040 27060 26160
rect 27180 26040 27300 26160
rect 27420 26040 27540 26160
rect 27660 26040 27780 26160
rect 27900 26040 28020 26160
rect 28140 26040 28260 26160
rect 28380 26040 28740 26160
rect 28860 26040 28980 26160
rect 29100 26040 29220 26160
rect 29340 26040 29460 26160
rect 29580 26040 29700 26160
rect 29820 26040 29940 26160
rect 30060 26040 30180 26160
rect 30300 26040 30420 26160
rect 30540 26040 30660 26160
rect 30780 26040 30900 26160
rect 31020 26040 31140 26160
rect 31260 26040 31380 26160
rect 31500 26040 31620 26160
rect 31740 26040 31860 26160
rect 31980 26040 32100 26160
rect 32220 26040 32580 26160
rect 32700 26040 32820 26160
rect 32940 26040 33060 26160
rect 33180 26040 33300 26160
rect 33420 26040 33540 26160
rect 33660 26040 33780 26160
rect 33900 26040 34020 26160
rect 34140 26040 34260 26160
rect 34380 26040 34500 26160
rect 34620 26040 34740 26160
rect 34860 26040 34980 26160
rect 35100 26040 35220 26160
rect 35340 26040 35460 26160
rect 35580 26040 35700 26160
rect 35820 26040 35940 26160
rect 36060 26040 36420 26160
rect 36540 26040 36660 26160
rect 36780 26040 36900 26160
rect 37020 26040 37140 26160
rect 37260 26040 37380 26160
rect 37500 26040 37620 26160
rect 37740 26040 37860 26160
rect 37980 26040 38100 26160
rect 38220 26040 38340 26160
rect 38460 26040 38580 26160
rect 38700 26040 38820 26160
rect 38940 26040 39060 26160
rect 39180 26040 39300 26160
rect 39420 26040 39540 26160
rect 39660 26040 39780 26160
rect 39900 26040 40020 26160
rect 40140 26040 40260 26160
rect 40380 26040 40500 26160
rect 40620 26040 40740 26160
rect 40860 26040 40980 26160
rect 41100 26040 41220 26160
rect 41340 26040 41460 26160
rect 41580 26040 41700 26160
rect 41820 26040 41940 26160
rect 42060 26040 42180 26160
rect 42300 26040 42420 26160
rect 42540 26040 42660 26160
rect 42780 26040 42900 26160
rect 43020 26040 43140 26160
rect 43260 26040 43380 26160
rect 43500 26040 43620 26160
rect 43740 26040 43860 26160
rect 43980 26040 44100 26160
rect 44220 26040 44340 26160
rect 44460 26040 44820 26160
rect 44940 26040 45060 26160
rect 45180 26040 45300 26160
rect 45420 26040 45540 26160
rect 45660 26040 45780 26160
rect 45900 26040 46020 26160
rect 46140 26040 46260 26160
rect 46380 26040 46500 26160
rect 46620 26040 46740 26160
rect 46860 26040 46980 26160
rect 47100 26040 47220 26160
rect 47340 26040 47460 26160
rect 47580 26040 47700 26160
rect 47820 26040 47940 26160
rect 48060 26040 48180 26160
rect 48300 26040 48420 26160
rect 48540 26040 48660 26160
rect 48780 26040 48900 26160
rect 49020 26040 49140 26160
rect 49260 26040 49380 26160
rect 49500 26040 49620 26160
rect 49740 26040 49860 26160
rect 49980 26040 50100 26160
rect 50220 26040 51330 26160
rect 52200 26040 52260 26160
rect 3135 26010 52260 26040
rect 5610 25920 5730 26010
rect 5340 25906 5460 25920
rect 5580 25876 5730 25920
rect 5580 25454 5594 25876
rect 5716 25454 5730 25876
rect 5580 25410 5730 25454
rect 6000 25860 6240 25920
rect 6000 25440 6060 25860
rect 6180 25440 6240 25860
rect 6000 25380 6240 25440
rect 6510 25876 6660 26010
rect 6510 25454 6524 25876
rect 6646 25454 6660 25876
rect 6510 25410 6660 25454
rect 6780 25906 6900 25920
rect 5340 25320 5460 25334
rect 5340 25230 5610 25320
rect 5340 24990 5460 25110
rect 6150 25080 6240 25380
rect 6780 25320 6900 25334
rect 7020 25906 7140 26010
rect 7410 25906 7530 25920
rect 7020 25320 7140 25334
rect 7260 25334 7410 25410
rect 7260 25320 7530 25334
rect 7740 25906 7860 25920
rect 7740 25320 7860 25334
rect 7980 25906 8100 25920
rect 8220 25890 8340 26010
rect 8220 25440 8340 25470
rect 8460 25906 8580 25920
rect 8100 25334 8460 25350
rect 7980 25320 8580 25334
rect 8700 25906 8820 26010
rect 9690 25920 9810 26010
rect 9090 25906 9210 25920
rect 8700 25320 8820 25334
rect 8940 25334 9090 25410
rect 8940 25320 9210 25334
rect 9420 25906 9540 25920
rect 9660 25876 9810 25920
rect 9660 25454 9674 25876
rect 9796 25454 9810 25876
rect 9660 25410 9810 25454
rect 10080 25860 10320 25920
rect 10080 25440 10140 25860
rect 10260 25440 10320 25860
rect 10080 25380 10320 25440
rect 10590 25876 10740 26010
rect 10590 25454 10604 25876
rect 10726 25454 10740 25876
rect 10590 25410 10740 25454
rect 10860 25906 10980 25920
rect 9420 25320 9540 25334
rect 6660 25230 6900 25320
rect 5580 25050 5670 25080
rect 5580 24960 5880 25050
rect 6090 24990 6240 25080
rect 6360 25110 6450 25170
rect 7020 24990 7140 25110
rect 6090 24810 6180 24990
rect 6060 24690 6180 24810
rect 6090 24480 6180 24690
rect 7260 24795 7380 25320
rect 7770 25110 7860 25320
rect 8010 25260 8550 25320
rect 7740 24990 8130 25110
rect 8340 25020 8460 25050
rect 8700 24990 8820 25110
rect 7260 24705 7845 24795
rect 5340 24466 5610 24480
rect 5460 24390 5610 24466
rect 6000 24466 6240 24480
rect 5340 23280 5460 23294
rect 5580 24210 5730 24270
rect 5580 23340 5594 24210
rect 5716 23340 5730 24210
rect 5580 23280 5730 23340
rect 6000 23294 6060 24466
rect 6180 23294 6240 24466
rect 6660 24466 6900 24480
rect 6660 24390 6780 24466
rect 6000 23280 6240 23294
rect 6510 24210 6660 24270
rect 6510 23340 6524 24210
rect 6646 23340 6660 24210
rect 5610 23190 5730 23280
rect 6510 23190 6660 23340
rect 6780 23280 6900 23294
rect 7020 23866 7140 23880
rect 7020 23190 7140 23294
rect 7260 23866 7380 24705
rect 7755 24510 7845 24705
rect 7500 24390 7620 24510
rect 7740 24480 7860 24510
rect 8040 24480 8130 24990
rect 8220 24795 8340 24810
rect 8715 24795 8805 24990
rect 8220 24705 8805 24795
rect 8220 24690 8340 24705
rect 8700 24495 8820 24510
rect 8940 24495 9060 25320
rect 9420 25230 9690 25320
rect 9300 25005 9420 25095
rect 10230 25080 10320 25380
rect 12060 25906 12180 26010
rect 12060 25620 12180 25634
rect 12300 25906 12420 25920
rect 10860 25320 10980 25334
rect 10740 25230 10980 25320
rect 12060 25290 12180 25410
rect 12300 25320 12420 25334
rect 12690 25906 12810 26010
rect 13980 25920 14100 26010
rect 12690 25320 12810 25334
rect 13020 25395 13140 25410
rect 13740 25395 13860 25650
rect 14940 25906 15060 25920
rect 13980 25620 14100 25650
rect 14715 25605 14940 25695
rect 9660 25050 9750 25080
rect 9660 24960 9960 25050
rect 10170 24990 10320 25080
rect 10440 25110 10530 25170
rect 10860 25095 10980 25110
rect 10860 25005 11925 25095
rect 10860 24990 10980 25005
rect 10170 24810 10260 24990
rect 10140 24690 10260 24810
rect 11835 24795 11925 25005
rect 12060 24795 12180 24810
rect 11835 24780 12180 24795
rect 12330 24780 12420 25320
rect 13020 25305 13860 25395
rect 13020 25290 13140 25305
rect 12540 25095 12660 25110
rect 13500 25095 13620 25110
rect 12540 25005 13620 25095
rect 12540 24990 12660 25005
rect 13500 24990 13620 25005
rect 12780 24795 12900 24810
rect 13500 24795 13620 24810
rect 12780 24780 13620 24795
rect 11835 24705 12420 24780
rect 12060 24690 12420 24705
rect 12660 24750 13620 24780
rect 7740 24390 7950 24480
rect 8040 24466 8190 24480
rect 8040 24390 8070 24466
rect 7860 24210 7950 24390
rect 7260 23280 7380 23294
rect 7500 23866 7620 23880
rect 7500 23190 7620 23294
rect 7830 23866 7950 23880
rect 7830 23190 7950 23294
rect 8070 23280 8190 23294
rect 8460 24466 8580 24480
rect 8700 24405 9060 24495
rect 8700 24390 8820 24405
rect 8460 23190 8580 23294
rect 8700 23866 8820 23880
rect 8700 23190 8820 23294
rect 8940 23866 9060 24405
rect 10170 24480 10260 24690
rect 12090 24480 12180 24690
rect 12780 24705 13620 24750
rect 12780 24690 12900 24705
rect 13500 24690 13620 24705
rect 9420 24466 9690 24480
rect 8940 23280 9060 23294
rect 9180 23866 9300 23880
rect 9180 23190 9300 23294
rect 9540 24390 9690 24466
rect 10080 24466 10320 24480
rect 9420 23280 9540 23294
rect 9660 24210 9810 24270
rect 9660 23340 9674 24210
rect 9796 23340 9810 24210
rect 9660 23280 9810 23340
rect 10080 23294 10140 24466
rect 10260 23294 10320 24466
rect 10740 24466 10980 24480
rect 10740 24390 10860 24466
rect 10080 23280 10320 23294
rect 10590 24210 10740 24270
rect 10590 23340 10604 24210
rect 10726 23340 10740 24210
rect 9690 23190 9810 23280
rect 10590 23190 10740 23340
rect 10860 23280 10980 23294
rect 12060 24466 12180 24480
rect 12060 23280 12180 23294
rect 12300 24466 12900 24480
rect 12420 24390 12900 24466
rect 12780 24346 12900 24390
rect 12300 23280 12420 23294
rect 12780 23280 12900 23324
rect 13740 23880 13860 25305
rect 13980 25395 14100 25410
rect 14715 25395 14805 25605
rect 13980 25305 14805 25395
rect 14940 25320 15060 25334
rect 15180 25906 15300 25920
rect 15420 25890 15540 26010
rect 15420 25440 15540 25470
rect 15660 25906 15780 25920
rect 15300 25334 15660 25350
rect 15180 25320 15780 25334
rect 20790 25906 20910 25920
rect 21180 25906 21300 26010
rect 20910 25334 21060 25410
rect 20790 25320 21060 25334
rect 21180 25320 21300 25334
rect 23100 25906 23220 26010
rect 23490 25906 23610 25920
rect 23100 25320 23220 25334
rect 13980 25290 14100 25305
rect 14970 25110 15060 25320
rect 15210 25260 15750 25320
rect 14940 24990 15330 25110
rect 15540 25020 15660 25050
rect 14940 24495 15060 24510
rect 14100 24480 15060 24495
rect 15240 24480 15330 24990
rect 14100 24405 15150 24480
rect 14940 24390 15150 24405
rect 15240 24466 15390 24480
rect 15240 24390 15270 24466
rect 15060 24210 15150 24390
rect 13740 23280 13860 23310
rect 12540 23190 12660 23280
rect 13980 23190 14100 23310
rect 15030 23866 15150 23880
rect 15030 23190 15150 23294
rect 15270 23280 15390 23294
rect 15660 24466 15780 24480
rect 18900 24405 19740 24495
rect 20700 24495 20820 24510
rect 19860 24405 20820 24495
rect 20700 24390 20820 24405
rect 20940 24495 21060 25320
rect 23460 25334 23490 25410
rect 23460 25320 23610 25334
rect 25500 25906 25620 25920
rect 25740 25876 25890 26010
rect 26670 25920 26790 26010
rect 25740 25454 25754 25876
rect 25876 25454 25890 25876
rect 25740 25410 25890 25454
rect 26160 25860 26400 25920
rect 26160 25440 26220 25860
rect 26340 25440 26400 25860
rect 25500 25320 25620 25334
rect 26160 25380 26400 25440
rect 26670 25876 26820 25920
rect 26670 25454 26684 25876
rect 26806 25454 26820 25876
rect 26670 25410 26820 25454
rect 26940 25906 27060 25920
rect 23100 25095 23220 25110
rect 22020 25005 23220 25095
rect 23100 24990 23220 25005
rect 23100 24495 23220 24510
rect 20940 24405 23220 24495
rect 15660 23190 15780 23294
rect 20700 23866 20820 23880
rect 20700 23190 20820 23294
rect 20940 23866 21060 24405
rect 23100 24390 23220 24405
rect 20940 23280 21060 23294
rect 21180 23866 21300 23880
rect 21180 23190 21300 23294
rect 23100 23866 23220 23880
rect 23100 23190 23220 23294
rect 23340 23866 23460 25290
rect 25500 25230 25740 25320
rect 25950 25110 26040 25170
rect 24300 25095 24420 25110
rect 25500 25095 25620 25110
rect 24300 25005 25620 25095
rect 24300 24990 24420 25005
rect 25500 24990 25620 25005
rect 26160 25080 26250 25380
rect 26940 25320 27060 25334
rect 27900 25906 28020 25920
rect 27900 25320 28020 25334
rect 28140 25906 28260 25920
rect 28380 25890 28500 26010
rect 30540 25920 30660 26010
rect 28380 25440 28500 25470
rect 28620 25906 28740 25920
rect 28260 25334 28620 25350
rect 28140 25320 28740 25334
rect 26790 25230 27060 25320
rect 27930 25110 28020 25320
rect 28170 25260 28710 25320
rect 26160 24990 26310 25080
rect 26730 25050 26820 25080
rect 26220 24810 26310 24990
rect 26520 24960 26820 25050
rect 26940 25095 27060 25110
rect 26940 25005 27420 25095
rect 26940 24990 27060 25005
rect 27900 25095 28290 25110
rect 27540 25005 28290 25095
rect 28620 25095 28740 25110
rect 28620 25050 29340 25095
rect 28500 25020 29340 25050
rect 27900 24990 28290 25005
rect 28620 25005 29340 25020
rect 28620 24990 28740 25005
rect 23700 24705 24540 24795
rect 26220 24690 26340 24810
rect 23580 24390 23700 24510
rect 26220 24480 26310 24690
rect 25500 24466 25740 24480
rect 23340 23280 23460 23294
rect 23580 23866 23700 23880
rect 23580 23190 23700 23294
rect 25620 24390 25740 24466
rect 26160 24466 26400 24480
rect 25500 23280 25620 23294
rect 25740 24210 25890 24270
rect 25740 23340 25754 24210
rect 25876 23340 25890 24210
rect 25740 23190 25890 23340
rect 26160 23294 26220 24466
rect 26340 23294 26400 24466
rect 26790 24466 27060 24480
rect 26790 24390 26940 24466
rect 26160 23280 26400 23294
rect 26670 24210 26820 24270
rect 26670 23340 26684 24210
rect 26806 23340 26820 24210
rect 26670 23280 26820 23340
rect 28200 24480 28290 24990
rect 28380 24795 28500 24810
rect 30300 24795 30420 25650
rect 30540 25620 30660 25650
rect 31020 25906 31140 25920
rect 30540 25290 30660 25410
rect 31020 25320 31140 25334
rect 31260 25906 31380 25920
rect 31500 25890 31620 26010
rect 32460 25920 32580 26010
rect 31500 25440 31620 25470
rect 31740 25906 31860 25920
rect 31380 25334 31740 25350
rect 31260 25320 31860 25334
rect 31050 25110 31140 25320
rect 31290 25260 31830 25320
rect 30540 25095 30660 25110
rect 31020 25095 31410 25110
rect 30540 25005 31410 25095
rect 31620 25020 31740 25050
rect 30540 24990 30660 25005
rect 31020 24990 31410 25005
rect 28380 24705 30420 24795
rect 28380 24690 28500 24705
rect 28020 24210 28110 24480
rect 28200 24466 28350 24480
rect 28200 24390 28230 24466
rect 26940 23280 27060 23294
rect 27990 23866 28110 23880
rect 26670 23190 26790 23280
rect 27990 23190 28110 23294
rect 28230 23280 28350 23294
rect 28620 24466 28740 24480
rect 28620 23190 28740 23294
rect 30300 23880 30420 24705
rect 30900 24405 31020 24495
rect 31320 24480 31410 24990
rect 31500 24795 31620 24810
rect 32220 24795 32340 25650
rect 32460 25620 32580 25650
rect 33180 25906 33300 26010
rect 33570 25906 33690 25920
rect 33180 25320 33300 25334
rect 33420 25334 33570 25410
rect 33420 25320 33690 25334
rect 34620 25906 34740 26010
rect 35010 25906 35130 25920
rect 34620 25320 34740 25334
rect 34860 25334 35010 25410
rect 36060 25906 36180 26010
rect 35130 25334 35820 25395
rect 33180 24990 33300 25110
rect 31500 24705 32340 24795
rect 31500 24690 31620 24705
rect 31140 24210 31230 24480
rect 31320 24466 31470 24480
rect 31320 24390 31350 24466
rect 30300 23280 30420 23310
rect 30540 23190 30660 23310
rect 31110 23866 31230 23880
rect 31110 23190 31230 23294
rect 31350 23280 31470 23294
rect 31740 24466 31860 24480
rect 31740 23190 31860 23294
rect 32220 23880 32340 24705
rect 33420 24795 33540 25320
rect 34860 25305 35820 25334
rect 32580 24705 33540 24795
rect 32220 23280 32340 23310
rect 32460 23190 32580 23310
rect 33180 23866 33300 23880
rect 33180 23190 33300 23294
rect 33420 23866 33540 24705
rect 33660 24495 33780 24510
rect 33660 24405 34620 24495
rect 33660 24390 33780 24405
rect 33420 23280 33540 23294
rect 33660 23866 33780 23880
rect 33660 23190 33780 23294
rect 34620 23866 34740 23880
rect 34620 23190 34740 23294
rect 34860 23866 34980 25305
rect 36450 25906 36570 25920
rect 36060 25320 36180 25334
rect 36300 25334 36450 25410
rect 36300 25320 36570 25334
rect 37500 25906 37620 26010
rect 37890 25906 38010 25920
rect 37500 25320 37620 25334
rect 37740 25334 37890 25410
rect 38940 25906 39060 26010
rect 38700 25395 38820 25410
rect 38010 25334 38820 25395
rect 34860 23280 34980 23294
rect 35100 23866 35220 23880
rect 35100 23190 35220 23294
rect 36060 23866 36180 23880
rect 36060 23190 36180 23294
rect 36300 23866 36420 25320
rect 37740 25305 38820 25334
rect 39330 25906 39450 25920
rect 38940 25320 39060 25334
rect 39180 25334 39330 25410
rect 40380 25906 40500 26010
rect 40140 25395 40260 25410
rect 39450 25334 40260 25395
rect 37500 25095 37620 25110
rect 36660 25005 37620 25095
rect 37500 24990 37620 25005
rect 36660 24405 36780 24495
rect 36300 23280 36420 23294
rect 36540 23866 36660 23880
rect 36540 23190 36660 23294
rect 37500 23866 37620 23880
rect 37500 23190 37620 23294
rect 37740 23866 37860 25305
rect 38700 25290 38820 25305
rect 39180 25305 40260 25334
rect 40770 25906 40890 25920
rect 40380 25320 40500 25334
rect 40620 25334 40770 25410
rect 40620 25320 40890 25334
rect 41820 25906 41940 26010
rect 42210 25906 42330 25920
rect 41820 25320 41940 25334
rect 42060 25334 42210 25410
rect 43260 25906 43380 26010
rect 43260 25620 43380 25634
rect 43500 25906 43620 25920
rect 43500 25620 43620 25634
rect 43740 25906 43860 26010
rect 43740 25620 43860 25634
rect 44460 25920 44580 26010
rect 48090 25920 48210 26010
rect 44460 25620 44580 25650
rect 44700 25876 44820 25920
rect 44700 25710 44820 25754
rect 42060 25320 42330 25334
rect 38940 24990 39060 25110
rect 37980 24390 38100 24510
rect 37740 23280 37860 23294
rect 37980 23866 38100 23880
rect 37980 23190 38100 23294
rect 38940 23866 39060 23880
rect 38940 23190 39060 23294
rect 39180 23866 39300 25305
rect 40140 25290 40260 25305
rect 39420 25095 39540 25110
rect 40380 25095 40500 25110
rect 39420 25005 40500 25095
rect 39420 24990 39540 25005
rect 40380 24990 40500 25005
rect 39180 23280 39300 23294
rect 39420 23866 39540 23880
rect 39420 23190 39540 23294
rect 40380 23866 40500 23880
rect 40380 23190 40500 23294
rect 40620 23866 40740 25320
rect 40860 25095 40980 25110
rect 41820 25095 41940 25110
rect 40860 25005 41940 25095
rect 40860 24990 40980 25005
rect 41820 24990 41940 25005
rect 40860 24390 40980 24510
rect 40620 23280 40740 23294
rect 40860 23866 40980 23880
rect 40860 23190 40980 23294
rect 41820 23866 41940 23880
rect 41820 23190 41940 23294
rect 42060 23866 42180 25320
rect 43260 25395 43380 25410
rect 42660 25305 43380 25395
rect 43260 25290 43380 25305
rect 43530 25110 43620 25620
rect 44460 25395 44580 25410
rect 44100 25305 44580 25395
rect 44460 25290 44580 25305
rect 43500 25095 43620 25110
rect 44460 25095 44580 25110
rect 43500 25005 44580 25095
rect 43500 24990 43620 25005
rect 44460 24990 44580 25005
rect 43530 24480 43620 24990
rect 42060 23280 42180 23294
rect 42300 23866 42420 23880
rect 42300 23190 42420 23294
rect 43500 24360 43650 24480
rect 43260 23190 43380 23310
rect 44700 23880 44820 25590
rect 47820 25906 47940 25920
rect 48060 25876 48210 25920
rect 48060 25454 48074 25876
rect 48196 25454 48210 25876
rect 48060 25410 48210 25454
rect 48480 25860 48720 25920
rect 48480 25440 48540 25860
rect 48660 25440 48720 25860
rect 48480 25380 48720 25440
rect 48990 25876 49140 26010
rect 48990 25454 49004 25876
rect 49126 25454 49140 25876
rect 48990 25410 49140 25454
rect 49260 25906 49380 25920
rect 47820 25320 47940 25334
rect 47820 25230 48090 25320
rect 48630 25080 48720 25380
rect 49260 25320 49380 25334
rect 49140 25230 49380 25320
rect 48060 25050 48150 25080
rect 48060 24960 48360 25050
rect 48570 24990 48720 25080
rect 48840 25110 48930 25170
rect 49260 25095 49380 25110
rect 49260 25005 49500 25095
rect 49260 24990 49380 25005
rect 48570 24810 48660 24990
rect 48540 24690 48660 24810
rect 48570 24480 48660 24690
rect 43650 23280 43770 23310
rect 44460 23190 44580 23310
rect 44700 23280 44820 23310
rect 47820 24466 48090 24480
rect 47940 24390 48090 24466
rect 48480 24466 48720 24480
rect 47820 23280 47940 23294
rect 48060 24210 48210 24270
rect 48060 23340 48074 24210
rect 48196 23340 48210 24210
rect 48060 23280 48210 23340
rect 48480 23294 48540 24466
rect 48660 23294 48720 24466
rect 49140 24466 49380 24480
rect 49140 24390 49260 24466
rect 48480 23280 48720 23294
rect 48990 24210 49140 24270
rect 48990 23340 49004 24210
rect 49126 23340 49140 24210
rect 48090 23190 48210 23280
rect 48990 23190 49140 23340
rect 49260 23280 49380 23294
rect 1155 23160 54240 23190
rect 1155 23040 1214 23160
rect 2086 23040 5220 23160
rect 5340 23040 5700 23160
rect 5820 23040 6180 23160
rect 6300 23040 6660 23160
rect 6780 23040 6900 23160
rect 7020 23040 7140 23160
rect 7260 23040 7380 23160
rect 7500 23040 7620 23160
rect 7740 23040 7860 23160
rect 7980 23040 8100 23160
rect 8220 23040 8580 23160
rect 8700 23040 8820 23160
rect 8940 23040 9060 23160
rect 9180 23040 9300 23160
rect 9420 23040 9540 23160
rect 9660 23040 9780 23160
rect 9900 23040 10020 23160
rect 10140 23040 10260 23160
rect 10380 23040 10500 23160
rect 10620 23040 10740 23160
rect 10860 23040 10980 23160
rect 11100 23040 11220 23160
rect 11340 23040 11460 23160
rect 11580 23040 11700 23160
rect 11820 23040 11940 23160
rect 12060 23040 12180 23160
rect 12300 23040 12420 23160
rect 12540 23040 12660 23160
rect 12780 23040 12900 23160
rect 13020 23040 13140 23160
rect 13260 23040 13380 23160
rect 13500 23040 13620 23160
rect 13740 23040 13860 23160
rect 13980 23040 14100 23160
rect 14220 23040 14340 23160
rect 14460 23040 14580 23160
rect 14700 23040 14820 23160
rect 14940 23040 15060 23160
rect 15180 23040 15300 23160
rect 15420 23040 15540 23160
rect 15660 23040 15780 23160
rect 15900 23040 16020 23160
rect 16140 23040 16260 23160
rect 16380 23040 16500 23160
rect 16620 23040 16740 23160
rect 16860 23040 16980 23160
rect 17100 23040 17220 23160
rect 17340 23040 17460 23160
rect 17580 23040 17700 23160
rect 17820 23040 17940 23160
rect 18060 23040 18180 23160
rect 18300 23040 18420 23160
rect 18540 23040 18660 23160
rect 18780 23040 18900 23160
rect 19020 23040 19140 23160
rect 19260 23040 19380 23160
rect 19500 23040 19620 23160
rect 19740 23040 19860 23160
rect 19980 23040 20100 23160
rect 20220 23040 20340 23160
rect 20460 23040 20580 23160
rect 20700 23040 20820 23160
rect 20940 23040 21060 23160
rect 21180 23040 21300 23160
rect 21420 23040 21540 23160
rect 21660 23040 21780 23160
rect 21900 23040 22020 23160
rect 22140 23040 22260 23160
rect 22380 23040 22500 23160
rect 22620 23040 22740 23160
rect 22860 23040 22980 23160
rect 23100 23040 23220 23160
rect 23340 23040 23460 23160
rect 23580 23040 23700 23160
rect 23820 23040 23940 23160
rect 24060 23040 24180 23160
rect 24300 23040 24420 23160
rect 24540 23040 24660 23160
rect 24780 23040 24900 23160
rect 25020 23040 25140 23160
rect 25260 23040 25380 23160
rect 25500 23040 25620 23160
rect 25740 23040 25860 23160
rect 25980 23040 26100 23160
rect 26220 23040 26580 23160
rect 26700 23040 27060 23160
rect 27180 23040 27300 23160
rect 27420 23040 27540 23160
rect 27660 23040 27780 23160
rect 27900 23040 28260 23160
rect 28380 23040 28740 23160
rect 28860 23040 28980 23160
rect 29100 23040 29220 23160
rect 29340 23040 29460 23160
rect 29580 23040 29700 23160
rect 29820 23040 29940 23160
rect 30060 23040 30180 23160
rect 30300 23040 30660 23160
rect 30780 23040 30900 23160
rect 31020 23040 31140 23160
rect 31260 23040 31380 23160
rect 31500 23040 31620 23160
rect 31740 23040 31860 23160
rect 31980 23040 32100 23160
rect 32220 23040 32340 23160
rect 32460 23040 32580 23160
rect 32700 23040 32820 23160
rect 32940 23040 33060 23160
rect 33180 23040 33540 23160
rect 33660 23040 33780 23160
rect 33900 23040 34020 23160
rect 34140 23040 34260 23160
rect 34380 23040 34500 23160
rect 34620 23040 34980 23160
rect 35100 23040 35220 23160
rect 35340 23040 35460 23160
rect 35580 23040 35700 23160
rect 35820 23040 35940 23160
rect 36060 23040 36180 23160
rect 36300 23040 36420 23160
rect 36540 23040 36660 23160
rect 36780 23040 36900 23160
rect 37020 23040 37140 23160
rect 37260 23040 37380 23160
rect 37500 23040 37620 23160
rect 37740 23040 37860 23160
rect 37980 23040 38100 23160
rect 38220 23040 38340 23160
rect 38460 23040 38580 23160
rect 38700 23040 38820 23160
rect 38940 23040 39300 23160
rect 39420 23040 39540 23160
rect 39660 23040 39780 23160
rect 39900 23040 40020 23160
rect 40140 23040 40260 23160
rect 40380 23040 40740 23160
rect 40860 23040 40980 23160
rect 41100 23040 41220 23160
rect 41340 23040 41460 23160
rect 41580 23040 41700 23160
rect 41820 23040 41940 23160
rect 42060 23040 42180 23160
rect 42300 23040 42420 23160
rect 42540 23040 42660 23160
rect 42780 23040 42900 23160
rect 43020 23040 43140 23160
rect 43260 23040 43620 23160
rect 43740 23040 43860 23160
rect 43980 23040 44100 23160
rect 44220 23040 44340 23160
rect 44460 23040 44580 23160
rect 44700 23040 44820 23160
rect 44940 23040 45060 23160
rect 45180 23040 45300 23160
rect 45420 23040 45540 23160
rect 45660 23040 45780 23160
rect 45900 23040 46020 23160
rect 46140 23040 46260 23160
rect 46380 23040 46500 23160
rect 46620 23040 46740 23160
rect 46860 23040 46980 23160
rect 47100 23040 47220 23160
rect 47340 23040 47460 23160
rect 47580 23040 47700 23160
rect 47820 23040 47940 23160
rect 48060 23040 48180 23160
rect 48300 23040 48420 23160
rect 48540 23040 48660 23160
rect 48780 23040 48900 23160
rect 49020 23040 49140 23160
rect 49260 23040 49380 23160
rect 49500 23040 49620 23160
rect 49740 23040 49860 23160
rect 49980 23040 50100 23160
rect 50220 23040 53310 23160
rect 54180 23040 54240 23160
rect 1155 23010 54240 23040
rect 5610 22920 5730 23010
rect 5340 22906 5460 22920
rect 5580 22860 5730 22920
rect 5580 21990 5594 22860
rect 5716 21990 5730 22860
rect 5580 21930 5730 21990
rect 6000 22906 6240 22920
rect 5460 21734 5610 21810
rect 5340 21720 5610 21734
rect 6000 21734 6060 22906
rect 6180 21734 6240 22906
rect 6510 22860 6660 23010
rect 6510 21990 6524 22860
rect 6646 21990 6660 22860
rect 6510 21930 6660 21990
rect 6780 22906 6900 22920
rect 6000 21720 6240 21734
rect 6660 21734 6780 21810
rect 8220 22906 8340 23010
rect 8220 22320 8340 22334
rect 8460 22906 8580 22920
rect 6660 21720 6900 21734
rect 6090 21510 6180 21720
rect 6060 21390 6180 21510
rect 5340 21090 5460 21210
rect 5580 21150 5880 21240
rect 6090 21210 6180 21390
rect 8460 21495 8580 22334
rect 8700 22906 8820 23010
rect 8700 22320 8820 22334
rect 9660 22906 9780 23010
rect 9660 22320 9780 22334
rect 9900 22906 10020 22920
rect 8700 21795 8820 21810
rect 9900 21795 10020 22334
rect 10140 22906 10260 23010
rect 10140 22320 10260 22334
rect 11190 22906 11310 23010
rect 11190 22320 11310 22334
rect 11430 22906 11550 22920
rect 8700 21705 10020 21795
rect 8700 21690 8820 21705
rect 8460 21405 9660 21495
rect 5580 21120 5670 21150
rect 6090 21120 6240 21210
rect 5340 20880 5610 20970
rect 5340 20866 5460 20880
rect 6150 20820 6240 21120
rect 7020 21195 7140 21210
rect 8220 21195 8340 21210
rect 7020 21105 8340 21195
rect 7020 21090 7140 21105
rect 8220 21090 8340 21105
rect 6360 21030 6450 21090
rect 6660 20880 6900 20970
rect 8460 20880 8580 21405
rect 9660 21195 9780 21210
rect 9060 21105 9780 21195
rect 9660 21090 9780 21105
rect 9900 20880 10020 21705
rect 11220 21810 11310 21990
rect 10380 21795 10500 21810
rect 11100 21795 11310 21810
rect 10380 21720 11310 21795
rect 11400 21734 11430 21810
rect 11400 21720 11550 21734
rect 11820 22906 11940 23010
rect 14490 22920 14610 23010
rect 11820 21720 11940 21734
rect 14220 22906 14340 22920
rect 14460 22860 14610 22920
rect 14460 21990 14474 22860
rect 14596 21990 14610 22860
rect 14460 21930 14610 21990
rect 14880 22906 15120 22920
rect 14340 21734 14490 21810
rect 14220 21720 14490 21734
rect 14880 21734 14940 22906
rect 15060 21734 15120 22906
rect 15390 22860 15540 23010
rect 15390 21990 15404 22860
rect 15526 21990 15540 22860
rect 15390 21930 15540 21990
rect 15660 22906 15780 22920
rect 14880 21720 15120 21734
rect 15540 21734 15660 21810
rect 15540 21720 15780 21734
rect 16860 22890 16980 22920
rect 17100 22890 17220 23010
rect 18060 22906 18180 23010
rect 18060 22320 18180 22334
rect 18300 22906 18420 22920
rect 10380 21705 11220 21720
rect 10380 21690 10500 21705
rect 11100 21690 11220 21705
rect 11400 21210 11490 21720
rect 14970 21510 15060 21720
rect 14940 21390 15060 21510
rect 11100 21195 11490 21210
rect 10500 21105 11490 21195
rect 11820 21195 11940 21210
rect 11820 21180 12300 21195
rect 11100 21090 11490 21105
rect 11700 21150 12300 21180
rect 11130 20880 11220 21090
rect 11820 21105 12300 21150
rect 11820 21090 11940 21105
rect 14460 21150 14760 21240
rect 14970 21210 15060 21390
rect 14460 21120 14550 21150
rect 14970 21120 15120 21210
rect 11370 20880 11910 20940
rect 14220 20880 14490 20970
rect 5340 20280 5460 20294
rect 5580 20746 5730 20790
rect 5580 20324 5594 20746
rect 5716 20324 5730 20746
rect 5580 20280 5730 20324
rect 6000 20760 6240 20820
rect 6780 20866 6900 20880
rect 6000 20340 6060 20760
rect 6180 20340 6240 20760
rect 6000 20280 6240 20340
rect 6510 20746 6660 20790
rect 6510 20324 6524 20746
rect 6646 20324 6660 20746
rect 5610 20190 5730 20280
rect 6510 20190 6660 20324
rect 6780 20280 6900 20294
rect 8220 20866 8340 20880
rect 8460 20866 8730 20880
rect 8460 20790 8610 20866
rect 8220 20190 8340 20294
rect 8610 20280 8730 20294
rect 9660 20866 9780 20880
rect 9900 20866 10170 20880
rect 9900 20790 10050 20866
rect 9660 20190 9780 20294
rect 10050 20280 10170 20294
rect 11100 20866 11220 20880
rect 11100 20280 11220 20294
rect 11340 20866 11940 20880
rect 11460 20850 11820 20866
rect 11340 20280 11460 20294
rect 11580 20730 11700 20760
rect 11580 20190 11700 20310
rect 11820 20280 11940 20294
rect 14220 20866 14340 20880
rect 15030 20820 15120 21120
rect 15240 21030 15330 21090
rect 15540 20880 15780 20970
rect 14220 20280 14340 20294
rect 14460 20746 14610 20790
rect 14460 20324 14474 20746
rect 14596 20324 14610 20746
rect 14460 20280 14610 20324
rect 14880 20760 15120 20820
rect 15660 20866 15780 20880
rect 14880 20340 14940 20760
rect 15060 20340 15120 20760
rect 14880 20280 15120 20340
rect 15390 20746 15540 20790
rect 15390 20324 15404 20746
rect 15526 20324 15540 20746
rect 14490 20190 14610 20280
rect 15390 20190 15540 20324
rect 15660 20280 15780 20294
rect 16860 20610 16980 22320
rect 18300 20910 18420 22334
rect 18540 22906 18660 23010
rect 18540 22320 18660 22334
rect 18780 22906 18900 22920
rect 19020 22860 19170 23010
rect 19950 22920 20070 23010
rect 19020 21990 19034 22860
rect 19156 21990 19170 22860
rect 19020 21930 19170 21990
rect 19440 22906 19680 22920
rect 18900 21734 19020 21810
rect 18780 21720 19020 21734
rect 19440 21734 19500 22906
rect 19620 21734 19680 22906
rect 19950 22860 20100 22920
rect 19950 21990 19964 22860
rect 20086 21990 20100 22860
rect 19950 21930 20100 21990
rect 20220 22906 20340 22920
rect 19440 21720 19680 21734
rect 20070 21734 20220 21810
rect 20070 21720 20340 21734
rect 20460 22906 20580 22920
rect 20700 22860 20850 23010
rect 21630 22920 21750 23010
rect 20700 21990 20714 22860
rect 20836 21990 20850 22860
rect 20700 21930 20850 21990
rect 21120 22906 21360 22920
rect 20580 21734 20700 21810
rect 20460 21720 20700 21734
rect 21120 21734 21180 22906
rect 21300 21734 21360 22906
rect 21630 22860 21780 22920
rect 21630 21990 21644 22860
rect 21766 21990 21780 22860
rect 21630 21930 21780 21990
rect 21900 22906 22020 22920
rect 21120 21720 21360 21734
rect 21750 21734 21900 21810
rect 22230 22906 22350 23010
rect 22230 22320 22350 22334
rect 22470 22906 22590 22920
rect 21750 21720 22020 21734
rect 19500 21510 19590 21720
rect 19500 21390 19620 21510
rect 21180 21510 21270 21720
rect 22260 21720 22350 21990
rect 22440 21734 22470 21810
rect 22440 21720 22590 21734
rect 22860 22906 22980 23010
rect 25020 22890 25140 23010
rect 25260 22890 25380 22920
rect 26310 22906 26430 23010
rect 26310 22320 26430 22334
rect 26550 22906 26670 22920
rect 22860 21720 22980 21734
rect 21180 21390 21300 21510
rect 19500 21210 19590 21390
rect 19230 21030 19320 21090
rect 19440 21120 19590 21210
rect 19800 21150 20100 21240
rect 21180 21210 21270 21390
rect 20010 21120 20100 21150
rect 17100 20895 17220 20910
rect 17100 20805 17820 20895
rect 17100 20790 17220 20805
rect 18060 20866 18180 20880
rect 16860 20446 16980 20490
rect 16860 20280 16980 20324
rect 17100 20550 17220 20580
rect 17100 20190 17220 20280
rect 18780 20880 19020 20970
rect 18420 20866 18570 20880
rect 18420 20790 18450 20866
rect 18060 20190 18180 20294
rect 18450 20280 18570 20294
rect 18780 20866 18900 20880
rect 19440 20820 19530 21120
rect 20910 21030 21000 21090
rect 21120 21120 21270 21210
rect 21480 21150 21780 21240
rect 22440 21210 22530 21720
rect 25260 21495 25380 22320
rect 26340 21810 26430 21990
rect 25500 21795 25620 21810
rect 25500 21705 25980 21795
rect 25500 21690 25620 21705
rect 26220 21795 26430 21810
rect 26100 21720 26430 21795
rect 26520 21734 26550 21810
rect 26520 21720 26670 21734
rect 26940 22906 27060 23010
rect 27990 22906 28110 23010
rect 27990 22320 28110 22334
rect 28230 22906 28350 22920
rect 28020 21810 28110 21990
rect 26940 21720 27060 21734
rect 27900 21720 28110 21810
rect 28200 21734 28230 21810
rect 28200 21720 28350 21734
rect 28620 22906 28740 23010
rect 29100 22906 29220 23010
rect 29100 22320 29220 22334
rect 29340 22906 29460 22920
rect 28620 21720 28740 21734
rect 28860 21795 28980 21810
rect 29340 21795 29460 22334
rect 29580 22906 29700 23010
rect 29580 22320 29700 22334
rect 30300 22906 30420 23010
rect 26100 21705 26340 21720
rect 26220 21690 26340 21705
rect 26220 21495 26340 21510
rect 25260 21405 26340 21495
rect 21690 21120 21780 21150
rect 20070 20880 20340 20970
rect 20220 20866 20340 20880
rect 18780 20280 18900 20294
rect 19020 20746 19170 20790
rect 19020 20324 19034 20746
rect 19156 20324 19170 20746
rect 19020 20190 19170 20324
rect 19440 20760 19680 20820
rect 19440 20340 19500 20760
rect 19620 20340 19680 20760
rect 19440 20280 19680 20340
rect 19950 20746 20100 20790
rect 19950 20324 19964 20746
rect 20086 20324 20100 20746
rect 19950 20280 20100 20324
rect 20220 20280 20340 20294
rect 20460 20880 20700 20970
rect 20460 20866 20580 20880
rect 21120 20820 21210 21120
rect 22140 21090 22380 21210
rect 22500 21090 22530 21210
rect 22860 21195 22980 21210
rect 22860 21180 23445 21195
rect 22740 21150 23445 21180
rect 21750 20880 22020 20970
rect 22170 20880 22260 21090
rect 22860 21105 23445 21150
rect 22860 21090 22980 21105
rect 22410 20880 22950 20940
rect 23355 20895 23445 21105
rect 21900 20866 22020 20880
rect 20460 20280 20580 20294
rect 20700 20746 20850 20790
rect 20700 20324 20714 20746
rect 20836 20324 20850 20746
rect 19950 20190 20070 20280
rect 20700 20190 20850 20324
rect 21120 20760 21360 20820
rect 21120 20340 21180 20760
rect 21300 20340 21360 20760
rect 21120 20280 21360 20340
rect 21630 20746 21780 20790
rect 21630 20324 21644 20746
rect 21766 20324 21780 20746
rect 21630 20280 21780 20324
rect 21900 20280 22020 20294
rect 22140 20866 22260 20880
rect 22140 20280 22260 20294
rect 22380 20866 22980 20880
rect 22500 20850 22860 20866
rect 22380 20280 22500 20294
rect 22620 20730 22740 20760
rect 21630 20190 21750 20280
rect 22620 20190 22740 20310
rect 23355 20805 24300 20895
rect 25020 20895 25140 20910
rect 24420 20805 25140 20895
rect 25020 20790 25140 20805
rect 22860 20280 22980 20294
rect 25020 20550 25140 20580
rect 25260 20550 25380 21405
rect 26220 21390 26340 21405
rect 26520 21210 26610 21720
rect 27900 21690 28020 21720
rect 26700 21390 26820 21510
rect 28200 21210 28290 21720
rect 28860 21705 29460 21795
rect 28860 21690 28980 21705
rect 28500 21405 29205 21495
rect 29115 21210 29205 21405
rect 26220 21090 26610 21210
rect 26940 21195 27060 21210
rect 26940 21180 27420 21195
rect 26820 21150 27420 21180
rect 26250 20880 26340 21090
rect 26940 21105 27420 21150
rect 26940 21090 27060 21105
rect 27900 21090 28140 21210
rect 28260 21090 28290 21210
rect 28620 21195 28740 21210
rect 28860 21195 28980 21210
rect 28620 21180 28980 21195
rect 28500 21150 28980 21180
rect 26490 20880 27030 20940
rect 27930 20880 28020 21090
rect 28620 21105 28980 21150
rect 28620 21090 28740 21105
rect 28860 21090 28980 21105
rect 29100 21090 29220 21210
rect 28170 20880 28710 20940
rect 29340 20880 29460 21705
rect 29580 21795 29700 21810
rect 29580 21705 29820 21795
rect 29580 21690 29700 21705
rect 30300 21720 30420 21734
rect 30690 22906 30810 22920
rect 30930 22906 31050 23010
rect 30930 22320 31050 22334
rect 31980 22906 32100 23010
rect 31980 22320 32100 22334
rect 32220 22906 32340 22920
rect 30930 21810 31020 21990
rect 30810 21734 30840 21810
rect 30690 21720 30840 21734
rect 30930 21795 31140 21810
rect 32220 21795 32340 22334
rect 32460 22906 32580 23010
rect 32460 22320 32580 22334
rect 33180 22906 33300 23010
rect 33180 22320 33300 22334
rect 33420 22906 33540 22920
rect 30930 21720 32340 21795
rect 30540 21495 30660 21510
rect 29700 21405 30660 21495
rect 30540 21390 30660 21405
rect 30750 21210 30840 21720
rect 31020 21705 32340 21720
rect 31020 21690 31140 21705
rect 29820 21195 29940 21210
rect 30300 21195 30420 21210
rect 29820 21180 30420 21195
rect 29820 21150 30540 21180
rect 29820 21105 30420 21150
rect 29820 21090 29940 21105
rect 30300 21090 30420 21105
rect 30750 21090 30780 21210
rect 30900 21090 31140 21210
rect 31980 21195 32100 21210
rect 31380 21105 32100 21195
rect 31980 21090 32100 21105
rect 30330 20880 30870 20940
rect 31020 20880 31110 21090
rect 32220 20880 32340 21705
rect 33180 21195 33300 21210
rect 33060 21105 33300 21195
rect 33180 21090 33300 21105
rect 33420 21195 33540 22334
rect 33660 22906 33780 23010
rect 33660 22320 33780 22334
rect 34620 22906 34740 23010
rect 34620 22320 34740 22334
rect 34860 22906 34980 22920
rect 33420 21105 34620 21195
rect 33420 20910 33540 21105
rect 26220 20866 26340 20880
rect 26220 20280 26340 20294
rect 26460 20866 27060 20880
rect 26580 20850 26940 20866
rect 26460 20280 26580 20294
rect 26700 20730 26820 20760
rect 25020 20190 25140 20280
rect 26700 20190 26820 20310
rect 26940 20280 27060 20294
rect 27900 20866 28020 20880
rect 27900 20280 28020 20294
rect 28140 20866 28740 20880
rect 28260 20850 28620 20866
rect 28140 20280 28260 20294
rect 28380 20730 28500 20760
rect 28380 20190 28500 20310
rect 28620 20280 28740 20294
rect 29100 20866 29220 20880
rect 29340 20866 29610 20880
rect 29340 20790 29490 20866
rect 29100 20190 29220 20294
rect 29490 20280 29610 20294
rect 30300 20866 30900 20880
rect 30420 20850 30780 20866
rect 30300 20280 30420 20294
rect 30540 20730 30660 20760
rect 30540 20190 30660 20310
rect 30780 20280 30900 20294
rect 31020 20866 31140 20880
rect 31020 20280 31140 20294
rect 31980 20866 32100 20880
rect 32220 20866 32490 20880
rect 32220 20790 32370 20866
rect 31980 20190 32100 20294
rect 32370 20280 32490 20294
rect 33180 20866 33300 20880
rect 34860 20910 34980 22334
rect 35100 22906 35220 23010
rect 35100 22320 35220 22334
rect 35820 22906 35940 23010
rect 35820 22320 35940 22334
rect 36060 22906 36180 22920
rect 36060 21495 36180 22334
rect 36300 22906 36420 23010
rect 37050 22920 37170 23010
rect 36300 22320 36420 22334
rect 36780 22906 36900 22920
rect 36300 21795 36420 21810
rect 36300 21705 36540 21795
rect 36300 21690 36420 21705
rect 37020 22860 37170 22920
rect 37020 21990 37034 22860
rect 37156 21990 37170 22860
rect 37020 21930 37170 21990
rect 37440 22906 37680 22920
rect 36900 21734 37050 21810
rect 36780 21720 37050 21734
rect 37440 21734 37500 22906
rect 37620 21734 37680 22906
rect 37950 22860 38100 23010
rect 37950 21990 37964 22860
rect 38086 21990 38100 22860
rect 37950 21930 38100 21990
rect 38220 22906 38340 22920
rect 37440 21720 37680 21734
rect 38100 21734 38220 21810
rect 39030 22906 39150 23010
rect 39030 22320 39150 22334
rect 39270 22906 39390 22920
rect 39060 21810 39150 21990
rect 38100 21720 38340 21734
rect 38940 21720 39150 21810
rect 39240 21734 39270 21810
rect 39240 21720 39390 21734
rect 39660 22906 39780 23010
rect 40380 22906 40500 23010
rect 40380 22320 40500 22334
rect 40620 22906 40740 22920
rect 39660 21720 39780 21734
rect 39900 21795 40020 21810
rect 40620 21795 40740 22334
rect 40860 22906 40980 23010
rect 40860 22320 40980 22334
rect 41670 22906 41790 23010
rect 41670 22320 41790 22334
rect 41910 22906 42030 22920
rect 36780 21495 36900 21510
rect 36060 21405 36900 21495
rect 35820 21195 35940 21210
rect 35460 21105 35940 21195
rect 35820 21090 35940 21105
rect 33540 20866 33690 20880
rect 33540 20790 33570 20866
rect 33180 20190 33300 20294
rect 33570 20280 33690 20294
rect 34620 20866 34740 20880
rect 36060 20880 36180 21405
rect 36780 21390 36900 21405
rect 37530 21510 37620 21720
rect 38940 21690 39060 21720
rect 37500 21390 37620 21510
rect 36780 21090 36900 21210
rect 37020 21150 37320 21240
rect 37530 21210 37620 21390
rect 39240 21210 39330 21720
rect 39900 21705 40740 21795
rect 39900 21690 40020 21705
rect 39420 21495 39540 21510
rect 39420 21405 40245 21495
rect 39420 21390 39540 21405
rect 37020 21120 37110 21150
rect 37530 21120 37680 21210
rect 36780 20880 37050 20970
rect 34980 20866 35130 20880
rect 34980 20790 35010 20866
rect 34620 20190 34740 20294
rect 35010 20280 35130 20294
rect 35820 20866 35940 20880
rect 36060 20866 36330 20880
rect 36060 20790 36210 20866
rect 35820 20190 35940 20294
rect 36210 20280 36330 20294
rect 36780 20866 36900 20880
rect 37590 20820 37680 21120
rect 38220 21195 38340 21210
rect 38940 21195 39330 21210
rect 38220 21105 39330 21195
rect 38220 21090 38340 21105
rect 38940 21090 39330 21105
rect 39540 21150 39660 21180
rect 37800 21030 37890 21090
rect 38100 20880 38340 20970
rect 38970 20880 39060 21090
rect 40155 21195 40245 21405
rect 40155 21105 40380 21195
rect 39210 20880 39750 20940
rect 40620 20880 40740 21705
rect 41700 21810 41790 21990
rect 40860 21795 40980 21810
rect 40860 21705 41100 21795
rect 40860 21690 40980 21705
rect 41580 21795 41790 21810
rect 41220 21720 41790 21795
rect 41880 21734 41910 21810
rect 41880 21720 42030 21734
rect 42300 22906 42420 23010
rect 42300 21720 42420 21734
rect 43260 22890 43380 23010
rect 44490 22920 44610 23010
rect 43650 22890 43770 22920
rect 43500 21720 43650 21840
rect 44220 22906 44340 22920
rect 44460 22860 44610 22920
rect 44460 21990 44474 22860
rect 44596 21990 44610 22860
rect 44460 21930 44610 21990
rect 44880 22906 45120 22920
rect 44340 21734 44490 21810
rect 44220 21720 44490 21734
rect 44880 21734 44940 22906
rect 45060 21734 45120 22906
rect 45390 22860 45540 23010
rect 45390 21990 45404 22860
rect 45526 21990 45540 22860
rect 45390 21930 45540 21990
rect 45660 22906 45780 22920
rect 44880 21720 45120 21734
rect 45540 21734 45660 21810
rect 45540 21720 45780 21734
rect 45900 22906 46020 22920
rect 46140 22860 46290 23010
rect 47070 22920 47190 23010
rect 46140 21990 46154 22860
rect 46276 21990 46290 22860
rect 46140 21930 46290 21990
rect 46560 22906 46800 22920
rect 46020 21734 46140 21810
rect 45900 21720 46140 21734
rect 46560 21734 46620 22906
rect 46740 21734 46800 22906
rect 47070 22860 47220 22920
rect 47070 21990 47084 22860
rect 47206 21990 47220 22860
rect 47070 21930 47220 21990
rect 47340 22906 47460 22920
rect 46560 21720 46800 21734
rect 47190 21734 47340 21810
rect 47580 22890 47700 23010
rect 49500 22920 49620 23010
rect 47820 22890 47940 22920
rect 47190 21720 47460 21734
rect 41220 21705 41700 21720
rect 41580 21690 41700 21705
rect 41880 21210 41970 21720
rect 42060 21390 42180 21510
rect 43530 21210 43620 21720
rect 43740 21390 43860 21510
rect 44970 21510 45060 21720
rect 44940 21390 45060 21510
rect 41580 21090 41970 21210
rect 42180 21150 42300 21180
rect 41610 20880 41700 21090
rect 42540 21195 42660 21210
rect 42540 21105 43500 21195
rect 42540 21090 42660 21105
rect 44220 21195 44340 21210
rect 43860 21105 44340 21195
rect 44220 21090 44340 21105
rect 44460 21150 44760 21240
rect 44970 21210 45060 21390
rect 46620 21510 46710 21720
rect 46620 21390 46740 21510
rect 46620 21210 46710 21390
rect 44460 21120 44550 21150
rect 44970 21120 45120 21210
rect 41850 20880 42390 20940
rect 42780 20895 42900 20910
rect 43260 20895 43380 20910
rect 36780 20280 36900 20294
rect 37020 20746 37170 20790
rect 37020 20324 37034 20746
rect 37156 20324 37170 20746
rect 37020 20280 37170 20324
rect 37440 20760 37680 20820
rect 38220 20866 38340 20880
rect 37440 20340 37500 20760
rect 37620 20340 37680 20760
rect 37440 20280 37680 20340
rect 37950 20746 38100 20790
rect 37950 20324 37964 20746
rect 38086 20324 38100 20746
rect 37050 20190 37170 20280
rect 37950 20190 38100 20324
rect 38220 20280 38340 20294
rect 38940 20866 39060 20880
rect 38940 20280 39060 20294
rect 39180 20866 39780 20880
rect 39300 20850 39660 20866
rect 39180 20280 39300 20294
rect 39420 20730 39540 20760
rect 39420 20190 39540 20310
rect 39660 20280 39780 20294
rect 40380 20866 40500 20880
rect 40620 20866 40890 20880
rect 40620 20790 40770 20866
rect 40380 20190 40500 20294
rect 40770 20280 40890 20294
rect 41580 20866 41700 20880
rect 41580 20280 41700 20294
rect 41820 20866 42420 20880
rect 41940 20850 42300 20866
rect 41820 20280 41940 20294
rect 42060 20730 42180 20760
rect 42060 20190 42180 20310
rect 42780 20805 43380 20895
rect 42780 20790 42900 20805
rect 43260 20790 43380 20805
rect 43530 20580 43620 21090
rect 44220 20880 44490 20970
rect 44220 20866 44340 20880
rect 42300 20280 42420 20294
rect 43260 20566 43380 20580
rect 43260 20190 43380 20294
rect 43500 20566 43620 20580
rect 43500 20280 43620 20294
rect 43740 20566 43860 20580
rect 43740 20190 43860 20294
rect 45030 20820 45120 21120
rect 45660 21090 45780 21210
rect 45240 21030 45330 21090
rect 46350 21030 46440 21090
rect 46560 21120 46710 21210
rect 46920 21150 47220 21240
rect 47130 21120 47220 21150
rect 45540 20880 45780 20970
rect 44220 20280 44340 20294
rect 44460 20746 44610 20790
rect 44460 20324 44474 20746
rect 44596 20324 44610 20746
rect 44460 20280 44610 20324
rect 44880 20760 45120 20820
rect 45660 20866 45780 20880
rect 44880 20340 44940 20760
rect 45060 20340 45120 20760
rect 44880 20280 45120 20340
rect 45390 20746 45540 20790
rect 45390 20324 45404 20746
rect 45526 20324 45540 20746
rect 44490 20190 44610 20280
rect 45390 20190 45540 20324
rect 45660 20280 45780 20294
rect 45900 20880 46140 20970
rect 45900 20866 46020 20880
rect 46560 20820 46650 21120
rect 47820 21195 47940 22320
rect 48780 22906 49380 22920
rect 48900 22830 49260 22906
rect 48780 21720 48900 21734
rect 49740 22876 49860 22920
rect 49740 21810 49860 21854
rect 49380 21734 49860 21810
rect 49260 21720 49860 21734
rect 49050 21630 49140 21720
rect 49050 21540 49350 21630
rect 48060 21495 48180 21510
rect 48780 21495 48900 21510
rect 48060 21405 48900 21495
rect 48060 21390 48180 21405
rect 48780 21390 48900 21405
rect 49260 21510 49350 21540
rect 49260 21390 49380 21510
rect 49740 21495 49860 21510
rect 49740 21450 49980 21495
rect 49620 21420 49980 21450
rect 49740 21405 49980 21420
rect 49740 21390 49860 21405
rect 49050 21210 49140 21270
rect 49020 21195 49140 21210
rect 47820 21105 49140 21195
rect 47190 20880 47460 20970
rect 47340 20866 47460 20880
rect 45900 20280 46020 20294
rect 46140 20746 46290 20790
rect 46140 20324 46154 20746
rect 46276 20324 46290 20746
rect 46140 20190 46290 20324
rect 46560 20760 46800 20820
rect 46560 20340 46620 20760
rect 46740 20340 46800 20760
rect 46560 20280 46800 20340
rect 47070 20746 47220 20790
rect 47070 20324 47084 20746
rect 47206 20324 47220 20746
rect 47070 20280 47220 20324
rect 47340 20280 47460 20294
rect 47580 20550 47700 20580
rect 47820 20550 47940 21105
rect 49020 21090 49140 21105
rect 49260 20880 49350 21390
rect 49500 21195 49620 21210
rect 49500 21105 49740 21195
rect 49500 21090 49620 21105
rect 48780 20866 48900 20880
rect 47070 20190 47190 20280
rect 47580 20190 47700 20280
rect 48780 20190 48900 20294
rect 49170 20866 49410 20880
rect 49170 20294 49230 20866
rect 49350 20294 49410 20866
rect 49170 20280 49410 20294
rect 49680 20866 49800 20880
rect 49680 20190 49800 20294
rect 3135 20160 52260 20190
rect 3135 20040 3194 20160
rect 4066 20040 5220 20160
rect 5340 20040 5460 20160
rect 5580 20040 5700 20160
rect 5820 20040 5940 20160
rect 6060 20040 6180 20160
rect 6300 20040 6420 20160
rect 6540 20040 6660 20160
rect 6780 20040 6900 20160
rect 7020 20040 7140 20160
rect 7260 20040 7380 20160
rect 7500 20040 7620 20160
rect 7740 20040 7860 20160
rect 7980 20040 8100 20160
rect 8220 20040 8340 20160
rect 8460 20040 8580 20160
rect 8700 20040 8820 20160
rect 8940 20040 9060 20160
rect 9180 20040 9300 20160
rect 9420 20040 9540 20160
rect 9660 20040 10020 20160
rect 10140 20040 10260 20160
rect 10380 20040 10500 20160
rect 10620 20040 10740 20160
rect 10860 20040 10980 20160
rect 11100 20040 11220 20160
rect 11340 20040 11460 20160
rect 11580 20040 11940 20160
rect 12060 20040 12180 20160
rect 12300 20040 12420 20160
rect 12540 20040 12660 20160
rect 12780 20040 12900 20160
rect 13020 20040 13140 20160
rect 13260 20040 13380 20160
rect 13500 20040 13620 20160
rect 13740 20040 13860 20160
rect 13980 20040 14100 20160
rect 14220 20040 14340 20160
rect 14460 20040 14580 20160
rect 14700 20040 14820 20160
rect 14940 20040 15060 20160
rect 15180 20040 15300 20160
rect 15420 20040 15540 20160
rect 15660 20040 15780 20160
rect 15900 20040 16020 20160
rect 16140 20040 16260 20160
rect 16380 20040 16500 20160
rect 16620 20040 16740 20160
rect 16860 20040 16980 20160
rect 17100 20040 17220 20160
rect 17340 20040 17460 20160
rect 17580 20040 17700 20160
rect 17820 20040 17940 20160
rect 18060 20040 18180 20160
rect 18300 20040 18420 20160
rect 18540 20040 18660 20160
rect 18780 20040 18900 20160
rect 19020 20040 19140 20160
rect 19260 20040 19380 20160
rect 19500 20040 19860 20160
rect 19980 20040 20100 20160
rect 20220 20040 20340 20160
rect 20460 20040 20580 20160
rect 20700 20040 20820 20160
rect 20940 20040 21060 20160
rect 21180 20040 21300 20160
rect 21420 20040 21540 20160
rect 21660 20040 21780 20160
rect 21900 20040 22020 20160
rect 22140 20040 22500 20160
rect 22620 20040 22740 20160
rect 22860 20040 22980 20160
rect 23100 20040 23220 20160
rect 23340 20040 23460 20160
rect 23580 20040 23700 20160
rect 23820 20040 23940 20160
rect 24060 20040 24180 20160
rect 24300 20040 24420 20160
rect 24540 20040 24660 20160
rect 24780 20040 24900 20160
rect 25020 20040 25380 20160
rect 25500 20040 25620 20160
rect 25740 20040 25860 20160
rect 25980 20040 26100 20160
rect 26220 20040 26580 20160
rect 26700 20040 27060 20160
rect 27180 20040 27300 20160
rect 27420 20040 27540 20160
rect 27660 20040 27780 20160
rect 27900 20040 28020 20160
rect 28140 20040 28260 20160
rect 28380 20040 28740 20160
rect 28860 20040 28980 20160
rect 29100 20040 29220 20160
rect 29340 20040 29460 20160
rect 29580 20040 29700 20160
rect 29820 20040 29940 20160
rect 30060 20040 30180 20160
rect 30300 20040 30420 20160
rect 30540 20040 30660 20160
rect 30780 20040 30900 20160
rect 31020 20040 31140 20160
rect 31260 20040 31380 20160
rect 31500 20040 31620 20160
rect 31740 20040 31860 20160
rect 31980 20040 32340 20160
rect 32460 20040 32580 20160
rect 32700 20040 32820 20160
rect 32940 20040 33060 20160
rect 33180 20040 33540 20160
rect 33660 20040 33780 20160
rect 33900 20040 34020 20160
rect 34140 20040 34260 20160
rect 34380 20040 34500 20160
rect 34620 20040 34740 20160
rect 34860 20040 34980 20160
rect 35100 20040 35220 20160
rect 35340 20040 35460 20160
rect 35580 20040 35700 20160
rect 35820 20040 36180 20160
rect 36300 20040 36420 20160
rect 36540 20040 36660 20160
rect 36780 20040 37140 20160
rect 37260 20040 37620 20160
rect 37740 20040 37860 20160
rect 37980 20040 38100 20160
rect 38220 20040 38340 20160
rect 38460 20040 38580 20160
rect 38700 20040 38820 20160
rect 38940 20040 39300 20160
rect 39420 20040 39540 20160
rect 39660 20040 39780 20160
rect 39900 20040 40020 20160
rect 40140 20040 40260 20160
rect 40380 20040 40740 20160
rect 40860 20040 40980 20160
rect 41100 20040 41220 20160
rect 41340 20040 41460 20160
rect 41580 20040 41940 20160
rect 42060 20040 42180 20160
rect 42300 20040 42420 20160
rect 42540 20040 42660 20160
rect 42780 20040 42900 20160
rect 43020 20040 43140 20160
rect 43260 20040 43620 20160
rect 43740 20040 43860 20160
rect 43980 20040 44100 20160
rect 44220 20040 44340 20160
rect 44460 20040 44580 20160
rect 44700 20040 44820 20160
rect 44940 20040 45060 20160
rect 45180 20040 45300 20160
rect 45420 20040 45540 20160
rect 45660 20040 45780 20160
rect 45900 20040 46020 20160
rect 46140 20040 46500 20160
rect 46620 20040 46740 20160
rect 46860 20040 46980 20160
rect 47100 20040 47220 20160
rect 47340 20040 47460 20160
rect 47580 20040 47940 20160
rect 48060 20040 48180 20160
rect 48300 20040 48420 20160
rect 48540 20040 48660 20160
rect 48780 20040 48900 20160
rect 49020 20040 49380 20160
rect 49500 20040 49860 20160
rect 49980 20040 50100 20160
rect 50220 20040 51330 20160
rect 52200 20040 52260 20160
rect 3135 20010 52260 20040
rect 5580 19906 5700 19920
rect 5460 19605 5580 19695
rect 5580 19320 5700 19334
rect 5820 19906 5940 19920
rect 6060 19890 6180 20010
rect 6060 19440 6180 19470
rect 6300 19906 6420 19920
rect 5940 19334 6300 19350
rect 5820 19320 6420 19334
rect 8940 19906 9060 19920
rect 9180 19876 9330 20010
rect 10110 19920 10230 20010
rect 11850 19920 11970 20010
rect 9180 19454 9194 19876
rect 9316 19454 9330 19876
rect 9180 19410 9330 19454
rect 9600 19860 9840 19920
rect 9600 19440 9660 19860
rect 9780 19440 9840 19860
rect 8940 19320 9060 19334
rect 9600 19380 9840 19440
rect 10110 19876 10260 19920
rect 10110 19454 10124 19876
rect 10246 19454 10260 19876
rect 10110 19410 10260 19454
rect 10380 19906 10500 19920
rect 5610 19110 5700 19320
rect 5850 19260 6390 19320
rect 8940 19230 9180 19320
rect 5580 18990 5970 19110
rect 9390 19110 9480 19170
rect 6300 19095 6420 19110
rect 6300 19050 6780 19095
rect 6180 19020 6780 19050
rect 6300 19005 6780 19020
rect 6300 18990 6420 19005
rect 9600 19080 9690 19380
rect 10380 19320 10500 19334
rect 10230 19230 10500 19320
rect 11580 19906 11700 19920
rect 11820 19876 11970 19920
rect 11820 19454 11834 19876
rect 11956 19454 11970 19876
rect 11820 19410 11970 19454
rect 12240 19860 12480 19920
rect 12240 19440 12300 19860
rect 12420 19440 12480 19860
rect 12240 19380 12480 19440
rect 12750 19876 12900 20010
rect 13770 19920 13890 20010
rect 12750 19454 12764 19876
rect 12886 19454 12900 19876
rect 12750 19410 12900 19454
rect 13020 19906 13140 19920
rect 11580 19320 11700 19334
rect 11580 19230 11790 19320
rect 12000 19170 12060 19260
rect 12000 19110 12090 19170
rect 9600 18990 9750 19080
rect 10170 19050 10260 19080
rect 5880 18480 5970 18990
rect 9660 18810 9750 18990
rect 9960 18960 10260 19050
rect 11580 19095 11700 19110
rect 11220 19005 11700 19095
rect 11580 18990 11700 19005
rect 11820 19020 12090 19110
rect 12180 18870 12270 18960
rect 9660 18690 9780 18810
rect 9660 18480 9750 18690
rect 12000 18780 12270 18870
rect 12390 18870 12480 19380
rect 13020 19320 13140 19334
rect 12900 19230 13140 19320
rect 13500 19906 13620 19920
rect 13740 19876 13890 19920
rect 13740 19454 13754 19876
rect 13876 19454 13890 19876
rect 13740 19410 13890 19454
rect 14160 19860 14400 19920
rect 14160 19440 14220 19860
rect 14340 19440 14400 19860
rect 14160 19380 14400 19440
rect 14670 19876 14820 20010
rect 14670 19454 14684 19876
rect 14806 19454 14820 19876
rect 14670 19410 14820 19454
rect 14940 19906 15060 19920
rect 13500 19320 13620 19334
rect 13500 19230 13770 19320
rect 12600 19110 12690 19170
rect 13020 19095 13140 19110
rect 13020 19005 13260 19095
rect 13020 18990 13140 19005
rect 14310 19080 14400 19380
rect 14940 19320 15060 19334
rect 15510 19906 15630 20010
rect 15510 19320 15630 19334
rect 15900 19906 16020 19920
rect 16140 19906 16260 20010
rect 16140 19620 16260 19634
rect 17820 19906 17940 19920
rect 15900 19320 16020 19334
rect 16140 19395 16260 19410
rect 14820 19230 15060 19320
rect 13740 19050 13830 19080
rect 13740 18960 14040 19050
rect 14250 18990 14400 19080
rect 14520 19110 14610 19170
rect 14940 19095 15060 19110
rect 15420 19095 15540 19110
rect 14940 19005 15540 19095
rect 14940 18990 15060 19005
rect 15420 18990 15540 19005
rect 12390 18810 12540 18870
rect 14250 18810 14340 18990
rect 15435 18810 15525 18990
rect 12390 18780 12660 18810
rect 12450 18690 12660 18780
rect 11820 18570 12210 18660
rect 11820 18480 11910 18570
rect 12450 18480 12540 18690
rect 14220 18690 14340 18810
rect 15420 18780 15540 18810
rect 15900 18780 15990 19320
rect 16140 19305 16860 19395
rect 16140 19290 16260 19305
rect 17820 19320 17940 19334
rect 18060 19906 18180 19920
rect 18300 19890 18420 20010
rect 18300 19440 18420 19470
rect 18540 19906 18660 19920
rect 18180 19334 18540 19350
rect 18060 19320 18660 19334
rect 19500 19906 19620 20010
rect 19890 19906 20010 19920
rect 19500 19320 19620 19334
rect 17850 19110 17940 19320
rect 18090 19260 18630 19320
rect 19860 19334 19890 19410
rect 19860 19320 20010 19334
rect 20940 19906 21060 20010
rect 21330 19906 21450 19920
rect 20940 19320 21060 19334
rect 21180 19334 21330 19410
rect 21180 19320 21450 19334
rect 22140 19906 22260 20010
rect 22530 19906 22650 19920
rect 22140 19320 22260 19334
rect 22380 19334 22530 19410
rect 23580 19906 23700 20010
rect 24810 19920 24930 20010
rect 22650 19334 23100 19395
rect 17820 18990 18210 19110
rect 18540 19050 18660 19110
rect 18420 19020 18660 19050
rect 18540 18990 18660 19020
rect 16140 18780 16260 18810
rect 15420 18750 15660 18780
rect 15420 18690 15540 18750
rect 14250 18480 14340 18690
rect 15900 18690 16260 18780
rect 16140 18480 16230 18690
rect 5700 18210 5790 18480
rect 5880 18466 6030 18480
rect 5880 18390 5910 18466
rect 5670 17866 5790 17880
rect 5670 17190 5790 17294
rect 5910 17280 6030 17294
rect 6300 18466 6420 18480
rect 6300 17190 6420 17294
rect 8940 18466 9180 18480
rect 9060 18390 9180 18466
rect 9600 18466 9840 18480
rect 8940 17280 9060 17294
rect 9180 18210 9330 18270
rect 9180 17340 9194 18210
rect 9316 17340 9330 18210
rect 9180 17190 9330 17340
rect 9600 17294 9660 18466
rect 9780 17294 9840 18466
rect 10230 18466 10500 18480
rect 10230 18390 10380 18466
rect 9600 17280 9840 17294
rect 10110 18210 10260 18270
rect 10110 17340 10124 18210
rect 10246 17340 10260 18210
rect 10110 17280 10260 17340
rect 10380 17280 10500 17294
rect 11580 18466 11790 18480
rect 11700 18390 11790 18466
rect 12240 18466 12540 18480
rect 11580 17280 11700 17294
rect 11820 18210 11970 18270
rect 11820 17340 11834 18210
rect 11956 17340 11970 18210
rect 11820 17280 11970 17340
rect 12240 17294 12300 18466
rect 12420 18390 12540 18466
rect 12420 17294 12480 18390
rect 12900 18466 13140 18480
rect 12900 18390 13020 18466
rect 12240 17280 12480 17294
rect 12750 18210 12900 18270
rect 12750 17340 12764 18210
rect 12886 17340 12900 18210
rect 10110 17190 10230 17280
rect 11850 17190 11970 17280
rect 12750 17190 12900 17340
rect 13020 17280 13140 17294
rect 13500 18466 13770 18480
rect 13620 18390 13770 18466
rect 14160 18466 14400 18480
rect 13500 17280 13620 17294
rect 13740 18210 13890 18270
rect 13740 17340 13754 18210
rect 13876 17340 13890 18210
rect 13740 17280 13890 17340
rect 14160 17294 14220 18466
rect 14340 17294 14400 18466
rect 14820 18466 15060 18480
rect 14820 18390 14940 18466
rect 14160 17280 14400 17294
rect 14670 18210 14820 18270
rect 14670 17340 14684 18210
rect 14806 17340 14820 18210
rect 13770 17190 13890 17280
rect 14670 17190 14820 17340
rect 14940 17280 15060 17294
rect 15420 18466 16020 18480
rect 15420 18390 15900 18466
rect 15420 18346 15540 18390
rect 15420 17280 15540 17324
rect 15900 17280 16020 17294
rect 16140 18466 16260 18480
rect 17820 18495 17940 18510
rect 16500 18480 17940 18495
rect 18120 18480 18210 18990
rect 18300 18690 18420 18810
rect 16500 18405 18030 18480
rect 17820 18390 18030 18405
rect 18120 18466 18270 18480
rect 18120 18390 18150 18466
rect 17940 18210 18030 18390
rect 16140 17280 16260 17294
rect 17910 17866 18030 17880
rect 15660 17190 15780 17280
rect 17910 17190 18030 17294
rect 18150 17280 18270 17294
rect 18540 18466 18660 18480
rect 18540 17190 18660 17294
rect 19500 17866 19620 17880
rect 19500 17190 19620 17294
rect 19740 17866 19860 19290
rect 19980 18495 20100 18510
rect 19980 18405 20220 18495
rect 19980 18390 20100 18405
rect 20940 18495 21060 18510
rect 20340 18405 21060 18495
rect 20940 18390 21060 18405
rect 21180 18195 21300 19320
rect 22380 19305 23100 19334
rect 22140 18990 22260 19110
rect 21420 18390 21540 18510
rect 20340 18105 21300 18195
rect 19740 17280 19860 17294
rect 19980 17866 20100 17880
rect 19980 17190 20100 17294
rect 20940 17866 21060 17880
rect 20940 17190 21060 17294
rect 21180 17866 21300 18105
rect 21180 17280 21300 17294
rect 21420 17866 21540 17880
rect 21420 17190 21540 17294
rect 22140 17866 22260 17880
rect 22140 17190 22260 17294
rect 22380 17866 22500 19305
rect 23970 19906 24090 19920
rect 23580 19320 23700 19334
rect 23820 19334 23970 19410
rect 23820 19320 24090 19334
rect 24540 19906 24660 19920
rect 24780 19876 24930 19920
rect 24780 19454 24794 19876
rect 24916 19454 24930 19876
rect 24780 19410 24930 19454
rect 25200 19860 25440 19920
rect 25200 19440 25260 19860
rect 25380 19440 25440 19860
rect 25200 19380 25440 19440
rect 25710 19876 25860 20010
rect 25710 19454 25724 19876
rect 25846 19454 25860 19876
rect 25710 19410 25860 19454
rect 25980 19906 26100 19920
rect 24540 19320 24660 19334
rect 22980 19005 23580 19095
rect 23820 19095 23940 19320
rect 24540 19230 24810 19320
rect 24300 19095 24420 19110
rect 23820 19005 24420 19095
rect 22620 18495 22740 18510
rect 23820 18495 23940 19005
rect 24300 18990 24420 19005
rect 25350 19080 25440 19380
rect 25980 19320 26100 19334
rect 26220 19906 26340 19920
rect 26460 19890 26580 20010
rect 27420 19920 27540 20010
rect 26460 19440 26580 19470
rect 26700 19906 26820 19920
rect 26340 19334 26700 19350
rect 26220 19320 26820 19334
rect 26940 19906 27060 19920
rect 26940 19320 27060 19334
rect 25860 19230 26100 19320
rect 26250 19260 26790 19320
rect 24780 19050 24870 19080
rect 24780 18960 25080 19050
rect 25290 18990 25440 19080
rect 25560 19110 25650 19170
rect 26220 19050 26340 19110
rect 26940 19110 27030 19320
rect 26220 19020 26460 19050
rect 26220 18990 26340 19020
rect 26670 18990 27060 19110
rect 25290 18810 25380 18990
rect 25260 18690 25380 18810
rect 26460 18690 26580 18810
rect 22620 18405 23940 18495
rect 22620 18390 22740 18405
rect 22380 17280 22500 17294
rect 22620 17866 22740 17880
rect 22620 17190 22740 17294
rect 23580 17866 23700 17880
rect 23580 17190 23700 17294
rect 23820 17866 23940 18405
rect 25290 18480 25380 18690
rect 26670 18480 26760 18990
rect 26940 18795 27060 18810
rect 27180 18795 27300 19650
rect 27420 19620 27540 19650
rect 28380 19906 28500 19920
rect 28380 19320 28500 19334
rect 28620 19906 28740 19920
rect 28860 19890 28980 20010
rect 28860 19440 28980 19470
rect 29100 19906 29220 19920
rect 28740 19334 29100 19350
rect 28620 19320 29220 19334
rect 30540 19906 30660 20010
rect 30930 19906 31050 19920
rect 30540 19320 30660 19334
rect 30780 19334 30930 19410
rect 30780 19320 31050 19334
rect 31980 19906 32100 20010
rect 32370 19906 32490 19920
rect 31980 19320 32100 19334
rect 32220 19334 32370 19410
rect 32220 19320 32490 19334
rect 33180 19906 33300 19920
rect 33420 19890 33540 20010
rect 33420 19440 33540 19470
rect 33660 19906 33780 19920
rect 33300 19334 33660 19350
rect 33180 19320 33780 19334
rect 33900 19906 34020 19920
rect 33900 19320 34020 19334
rect 35820 19906 35940 20010
rect 36210 19906 36330 19920
rect 35820 19320 35940 19334
rect 36060 19334 36210 19410
rect 36780 19906 36900 20010
rect 36780 19620 36900 19634
rect 37020 19906 37140 19920
rect 36060 19320 36330 19334
rect 36540 19395 36660 19410
rect 36780 19395 36900 19410
rect 28410 19110 28500 19320
rect 28650 19260 29190 19320
rect 28380 18990 28770 19110
rect 29100 19095 29220 19110
rect 29580 19095 29700 19110
rect 29100 19050 29700 19095
rect 28980 19020 29700 19050
rect 29100 19005 29700 19020
rect 29100 18990 29220 19005
rect 29580 18990 29700 19005
rect 29835 19005 30540 19095
rect 26940 18705 27300 18795
rect 26940 18690 27060 18705
rect 24540 18466 24810 18480
rect 23820 17280 23940 17294
rect 24060 17866 24180 17880
rect 24060 17190 24180 17294
rect 24660 18390 24810 18466
rect 25200 18466 25440 18480
rect 24540 17280 24660 17294
rect 24780 18210 24930 18270
rect 24780 17340 24794 18210
rect 24916 17340 24930 18210
rect 24780 17280 24930 17340
rect 25200 17294 25260 18466
rect 25380 17294 25440 18466
rect 25860 18466 26100 18480
rect 25860 18390 25980 18466
rect 25200 17280 25440 17294
rect 25710 18210 25860 18270
rect 25710 17340 25724 18210
rect 25846 17340 25860 18210
rect 24810 17190 24930 17280
rect 25710 17190 25860 17340
rect 25980 17280 26100 17294
rect 26220 18466 26340 18480
rect 26220 17190 26340 17294
rect 26610 18466 26760 18480
rect 26730 18390 26760 18466
rect 26850 18210 26940 18480
rect 27180 17880 27300 18705
rect 28380 18480 28500 18510
rect 28680 18480 28770 18990
rect 28860 18795 28980 18810
rect 29835 18795 29925 19005
rect 28860 18705 29925 18795
rect 28860 18690 28980 18705
rect 29340 18495 29460 18510
rect 30780 18495 30900 19320
rect 31020 19095 31140 19110
rect 31980 19095 32100 19110
rect 31020 19005 32100 19095
rect 31020 18990 31140 19005
rect 31980 18990 32100 19005
rect 32220 19095 32340 19320
rect 33210 19260 33750 19320
rect 32220 19005 32460 19095
rect 28380 18390 28590 18480
rect 28680 18466 28830 18480
rect 28680 18390 28710 18466
rect 28500 18210 28590 18390
rect 26610 17280 26730 17294
rect 26850 17866 26970 17880
rect 26850 17190 26970 17294
rect 27180 17280 27300 17310
rect 27420 17190 27540 17310
rect 28470 17866 28590 17880
rect 28470 17190 28590 17294
rect 28710 17280 28830 17294
rect 29100 18466 29220 18480
rect 29340 18405 30900 18495
rect 29340 18390 29460 18405
rect 29100 17190 29220 17294
rect 30540 17866 30660 17880
rect 30540 17190 30660 17294
rect 30780 17866 30900 18405
rect 30780 17280 30900 17294
rect 31020 17866 31140 17880
rect 31020 17190 31140 17294
rect 31980 17866 32100 17880
rect 31980 17190 32100 17294
rect 32220 17866 32340 19005
rect 33900 19110 33990 19320
rect 33300 19020 33420 19050
rect 33630 19095 34020 19110
rect 33630 19005 35580 19095
rect 33630 18990 34020 19005
rect 32460 18495 32580 18510
rect 32460 18405 32700 18495
rect 32460 18390 32580 18405
rect 33630 18480 33720 18990
rect 33900 18495 34020 18510
rect 33900 18480 34860 18495
rect 33180 18466 33300 18480
rect 32220 17280 32340 17294
rect 32460 17866 32580 17880
rect 32460 17190 32580 17294
rect 33180 17190 33300 17294
rect 33570 18466 33720 18480
rect 33690 18390 33720 18466
rect 33810 18405 34860 18480
rect 33810 18390 34020 18405
rect 33810 18210 33900 18390
rect 33570 17280 33690 17294
rect 33810 17866 33930 17880
rect 33810 17190 33930 17294
rect 35820 17866 35940 17880
rect 35820 17190 35940 17294
rect 36060 17866 36180 19320
rect 36540 19305 36900 19395
rect 37020 19320 37140 19334
rect 37410 19906 37530 20010
rect 37410 19320 37530 19334
rect 37980 19906 38100 20010
rect 38370 19906 38490 19920
rect 37980 19320 38100 19334
rect 38220 19334 38370 19410
rect 38220 19320 38490 19334
rect 38940 19906 39060 20010
rect 39330 19906 39450 19920
rect 38940 19320 39060 19334
rect 39180 19334 39330 19410
rect 40380 19906 40500 20010
rect 41580 19920 41700 20010
rect 39660 19395 39780 19410
rect 39450 19334 39780 19395
rect 36540 19290 36660 19305
rect 36780 19290 36900 19305
rect 36780 18780 36900 18810
rect 37050 18780 37140 19320
rect 36780 18690 37140 18780
rect 37380 18750 37500 18780
rect 36810 18480 36900 18690
rect 36780 18466 36900 18480
rect 36060 17280 36180 17294
rect 36300 17866 36420 17880
rect 36300 17190 36420 17294
rect 36780 17280 36900 17294
rect 37020 18466 37620 18480
rect 37140 18390 37620 18466
rect 37500 18346 37620 18390
rect 37020 17280 37140 17294
rect 38220 18195 38340 19320
rect 39180 19305 39780 19334
rect 40770 19906 40890 19920
rect 40380 19320 40500 19334
rect 38940 18990 39060 19110
rect 38460 18390 38580 18510
rect 37860 18105 38340 18195
rect 37500 17280 37620 17324
rect 37980 17866 38100 17880
rect 37260 17190 37380 17280
rect 37980 17190 38100 17294
rect 38220 17866 38340 18105
rect 38220 17280 38340 17294
rect 38460 17866 38580 17880
rect 38460 17190 38580 17294
rect 38940 17866 39060 17880
rect 38940 17190 39060 17294
rect 39180 17866 39300 19305
rect 39660 19290 39780 19305
rect 40740 19334 40770 19410
rect 41580 19620 41700 19650
rect 40740 19320 40890 19334
rect 41100 19395 41220 19410
rect 41580 19395 41700 19410
rect 41100 19305 41700 19395
rect 41100 19290 41220 19305
rect 41580 19290 41700 19305
rect 39420 19095 39540 19110
rect 39420 19005 40380 19095
rect 39420 18990 39540 19005
rect 39540 18405 39900 18495
rect 39180 17280 39300 17294
rect 39420 17866 39540 17880
rect 39420 17190 39540 17294
rect 40380 17866 40500 17880
rect 40380 17190 40500 17294
rect 40620 17866 40740 19290
rect 41820 17880 41940 19650
rect 42840 19906 42960 20010
rect 42840 19320 42960 19334
rect 43230 19906 43470 19920
rect 43230 19334 43290 19906
rect 43410 19334 43470 19906
rect 43230 19320 43470 19334
rect 43740 19906 43860 20010
rect 43740 19320 43860 19334
rect 44460 19906 44580 19920
rect 44700 19890 44820 20010
rect 44700 19440 44820 19470
rect 44940 19906 45060 19920
rect 44580 19334 44940 19350
rect 44460 19320 45060 19334
rect 45180 19906 45300 19920
rect 46140 19906 46260 20010
rect 45300 19605 45900 19695
rect 45180 19320 45300 19334
rect 46530 19906 46650 19920
rect 46140 19320 46260 19334
rect 46380 19334 46530 19410
rect 47580 19906 47700 20010
rect 47580 19620 47700 19634
rect 47820 19906 47940 19920
rect 47820 19620 47940 19634
rect 48060 19906 48180 20010
rect 48060 19620 48180 19634
rect 49020 19906 49140 19920
rect 46380 19320 46650 19334
rect 43020 19095 43140 19110
rect 42180 19005 43140 19095
rect 43020 18990 43140 19005
rect 43290 18810 43380 19320
rect 44490 19260 45030 19320
rect 43500 18990 43620 19110
rect 44100 19005 44460 19095
rect 45180 19110 45270 19320
rect 44580 19020 44700 19050
rect 44910 18990 45300 19110
rect 45420 19095 45540 19110
rect 46140 19095 46260 19110
rect 45420 19005 46260 19095
rect 45420 18990 45540 19005
rect 46140 18990 46260 19005
rect 43500 18930 43590 18990
rect 42780 18795 42900 18810
rect 42420 18780 42900 18795
rect 42420 18750 43020 18780
rect 42420 18705 42900 18750
rect 42780 18690 42900 18705
rect 43260 18690 43380 18810
rect 43290 18660 43380 18690
rect 43290 18570 43590 18660
rect 43500 18480 43590 18570
rect 44910 18480 45000 18990
rect 45180 18495 45300 18510
rect 46380 18495 46500 19320
rect 47580 19290 47700 19410
rect 47850 19110 47940 19620
rect 49260 19890 49380 20010
rect 49260 19440 49380 19470
rect 49500 19906 49620 19920
rect 49140 19334 49500 19350
rect 49020 19320 49620 19334
rect 49740 19906 49860 19920
rect 49740 19320 49860 19334
rect 49050 19260 49590 19320
rect 47820 19095 47940 19110
rect 47460 19005 47940 19095
rect 47820 18990 47940 19005
rect 49020 19095 49140 19110
rect 48180 19050 49140 19095
rect 49740 19110 49830 19320
rect 48180 19020 49260 19050
rect 48180 19005 49140 19020
rect 49020 18990 49140 19005
rect 49470 18990 49860 19110
rect 45180 18480 46500 18495
rect 40620 17280 40740 17294
rect 40860 17866 40980 17880
rect 40860 17190 40980 17294
rect 41580 17190 41700 17310
rect 41820 17280 41940 17310
rect 42780 18466 43380 18480
rect 42780 18390 43260 18466
rect 42780 18346 42900 18390
rect 42780 17280 42900 17324
rect 43740 18466 43860 18480
rect 43380 17294 43740 17370
rect 43260 17280 43860 17294
rect 44460 18466 44580 18480
rect 43020 17190 43140 17280
rect 44460 17190 44580 17294
rect 44850 18466 45000 18480
rect 44970 18390 45000 18466
rect 45090 18405 46500 18480
rect 45090 18390 45300 18405
rect 45090 18210 45180 18390
rect 44850 17280 44970 17294
rect 45090 17866 45210 17880
rect 45090 17190 45210 17294
rect 46140 17866 46260 17880
rect 46140 17190 46260 17294
rect 46380 17866 46500 18405
rect 46620 18390 46740 18510
rect 47850 18480 47940 18990
rect 48180 18705 49260 18795
rect 49470 18480 49560 18990
rect 49740 18480 49860 18510
rect 46380 17280 46500 17294
rect 46620 17866 46740 17880
rect 46620 17190 46740 17294
rect 47820 18360 47970 18480
rect 47580 17190 47700 17310
rect 47970 17280 48090 17310
rect 49020 18466 49140 18480
rect 49020 17190 49140 17294
rect 49410 18466 49560 18480
rect 49530 18390 49560 18466
rect 49650 18390 49860 18480
rect 49650 18210 49740 18390
rect 49410 17280 49530 17294
rect 49650 17866 49770 17880
rect 49650 17190 49770 17294
rect 1155 17160 54240 17190
rect 1155 17040 1214 17160
rect 2086 17040 5220 17160
rect 5340 17040 5460 17160
rect 5580 17040 5700 17160
rect 5820 17040 5940 17160
rect 6060 17040 6180 17160
rect 6300 17040 6420 17160
rect 6540 17040 6660 17160
rect 6780 17040 6900 17160
rect 7020 17040 7140 17160
rect 7260 17040 7380 17160
rect 7500 17040 7620 17160
rect 7740 17040 7860 17160
rect 7980 17040 8100 17160
rect 8220 17040 8340 17160
rect 8460 17040 8580 17160
rect 8700 17040 8820 17160
rect 8940 17040 9060 17160
rect 9180 17040 9300 17160
rect 9420 17040 9540 17160
rect 9660 17040 9780 17160
rect 9900 17040 10020 17160
rect 10140 17040 10260 17160
rect 10380 17040 10500 17160
rect 10620 17040 10740 17160
rect 10860 17040 10980 17160
rect 11100 17040 11220 17160
rect 11340 17040 11460 17160
rect 11580 17040 11940 17160
rect 12060 17040 12420 17160
rect 12540 17040 12660 17160
rect 12780 17040 12900 17160
rect 13020 17040 13140 17160
rect 13260 17040 13380 17160
rect 13500 17040 13620 17160
rect 13740 17040 13860 17160
rect 13980 17040 14100 17160
rect 14220 17040 14340 17160
rect 14460 17040 14580 17160
rect 14700 17040 14820 17160
rect 14940 17040 15060 17160
rect 15180 17040 15300 17160
rect 15420 17040 15780 17160
rect 15900 17040 16260 17160
rect 16380 17040 16500 17160
rect 16620 17040 16740 17160
rect 16860 17040 16980 17160
rect 17100 17040 17220 17160
rect 17340 17040 17460 17160
rect 17580 17040 17700 17160
rect 17820 17040 17940 17160
rect 18060 17040 18180 17160
rect 18300 17040 18420 17160
rect 18540 17040 18660 17160
rect 18780 17040 18900 17160
rect 19020 17040 19140 17160
rect 19260 17040 19380 17160
rect 19500 17040 19620 17160
rect 19740 17040 19860 17160
rect 19980 17040 20100 17160
rect 20220 17040 20340 17160
rect 20460 17040 20580 17160
rect 20700 17040 20820 17160
rect 20940 17040 21060 17160
rect 21180 17040 21300 17160
rect 21420 17040 21540 17160
rect 21660 17040 21780 17160
rect 21900 17040 22020 17160
rect 22140 17040 22500 17160
rect 22620 17040 22740 17160
rect 22860 17040 22980 17160
rect 23100 17040 23220 17160
rect 23340 17040 23460 17160
rect 23580 17040 23940 17160
rect 24060 17040 24180 17160
rect 24300 17040 24420 17160
rect 24540 17040 24660 17160
rect 24780 17040 24900 17160
rect 25020 17040 25380 17160
rect 25500 17040 25620 17160
rect 25740 17040 25860 17160
rect 25980 17040 26100 17160
rect 26220 17040 26340 17160
rect 26460 17040 26580 17160
rect 26700 17040 26820 17160
rect 26940 17040 27300 17160
rect 27420 17040 27540 17160
rect 27660 17040 27780 17160
rect 27900 17040 28020 17160
rect 28140 17040 28260 17160
rect 28380 17040 28500 17160
rect 28620 17040 28740 17160
rect 28860 17040 28980 17160
rect 29100 17040 29220 17160
rect 29340 17040 29460 17160
rect 29580 17040 29700 17160
rect 29820 17040 29940 17160
rect 30060 17040 30180 17160
rect 30300 17040 30420 17160
rect 30540 17040 30900 17160
rect 31020 17040 31140 17160
rect 31260 17040 31380 17160
rect 31500 17040 31620 17160
rect 31740 17040 31860 17160
rect 31980 17040 32100 17160
rect 32220 17040 32340 17160
rect 32460 17040 32580 17160
rect 32700 17040 32820 17160
rect 32940 17040 33060 17160
rect 33180 17040 33540 17160
rect 33660 17040 33780 17160
rect 33900 17040 34020 17160
rect 34140 17040 34260 17160
rect 34380 17040 34500 17160
rect 34620 17040 34740 17160
rect 34860 17040 34980 17160
rect 35100 17040 35220 17160
rect 35340 17040 35460 17160
rect 35580 17040 35700 17160
rect 35820 17040 35940 17160
rect 36060 17040 36180 17160
rect 36300 17040 36420 17160
rect 36540 17040 36660 17160
rect 36780 17040 36900 17160
rect 37020 17040 37140 17160
rect 37260 17040 37380 17160
rect 37500 17040 37620 17160
rect 37740 17040 37860 17160
rect 37980 17040 38100 17160
rect 38220 17040 38340 17160
rect 38460 17040 38580 17160
rect 38700 17040 38820 17160
rect 38940 17040 39300 17160
rect 39420 17040 39540 17160
rect 39660 17040 39780 17160
rect 39900 17040 40020 17160
rect 40140 17040 40260 17160
rect 40380 17040 40500 17160
rect 40620 17040 40740 17160
rect 40860 17040 40980 17160
rect 41100 17040 41220 17160
rect 41340 17040 41460 17160
rect 41580 17040 41940 17160
rect 42060 17040 42180 17160
rect 42300 17040 42420 17160
rect 42540 17040 42660 17160
rect 42780 17040 42900 17160
rect 43020 17040 43140 17160
rect 43260 17040 43380 17160
rect 43500 17040 43620 17160
rect 43740 17040 43860 17160
rect 43980 17040 44100 17160
rect 44220 17040 44340 17160
rect 44460 17040 44820 17160
rect 44940 17040 45300 17160
rect 45420 17040 45540 17160
rect 45660 17040 45780 17160
rect 45900 17040 46020 17160
rect 46140 17040 46500 17160
rect 46620 17040 46740 17160
rect 46860 17040 46980 17160
rect 47100 17040 47220 17160
rect 47340 17040 47460 17160
rect 47580 17040 47700 17160
rect 47820 17040 47940 17160
rect 48060 17040 48180 17160
rect 48300 17040 48420 17160
rect 48540 17040 48660 17160
rect 48780 17040 48900 17160
rect 49020 17040 49380 17160
rect 49500 17040 49860 17160
rect 49980 17040 50100 17160
rect 50220 17040 53310 17160
rect 54180 17040 54240 17160
rect 1155 17010 54240 17040
rect 6300 16906 6420 17010
rect 6300 16320 6420 16334
rect 6540 16906 6660 16920
rect 6060 15195 6180 15210
rect 6300 15195 6420 15210
rect 6060 15105 6420 15195
rect 6060 15090 6180 15105
rect 6300 15090 6420 15105
rect 6540 14910 6660 16334
rect 6780 16906 6900 17010
rect 8010 16920 8130 17010
rect 6780 16320 6900 16334
rect 7740 16906 7860 16920
rect 6780 15690 6900 15810
rect 7980 16860 8130 16920
rect 7980 15990 7994 16860
rect 8116 15990 8130 16860
rect 7980 15930 8130 15990
rect 8400 16906 8640 16920
rect 7860 15734 8010 15810
rect 7740 15720 8010 15734
rect 8400 15734 8460 16906
rect 8580 15734 8640 16906
rect 8910 16860 9060 17010
rect 9690 16920 9810 17010
rect 8910 15990 8924 16860
rect 9046 15990 9060 16860
rect 8910 15930 9060 15990
rect 9180 16906 9300 16920
rect 8400 15720 8640 15734
rect 9060 15734 9180 15810
rect 9060 15720 9300 15734
rect 9420 16906 9540 16920
rect 9660 16860 9810 16920
rect 9660 15990 9674 16860
rect 9796 15990 9810 16860
rect 9660 15930 9810 15990
rect 10080 16906 10320 16920
rect 9540 15734 9690 15810
rect 9420 15720 9690 15734
rect 10080 15734 10140 16906
rect 10260 15734 10320 16906
rect 10590 16860 10740 17010
rect 11370 16920 11490 17010
rect 10590 15990 10604 16860
rect 10726 15990 10740 16860
rect 10590 15930 10740 15990
rect 10860 16906 10980 16920
rect 10080 15720 10320 15734
rect 10740 15734 10860 15810
rect 10740 15720 10980 15734
rect 11100 16906 11220 16920
rect 11340 16860 11490 16920
rect 11340 15990 11354 16860
rect 11476 15990 11490 16860
rect 11340 15930 11490 15990
rect 11760 16906 12000 16920
rect 11220 15734 11310 15810
rect 11100 15720 11310 15734
rect 11760 15734 11820 16906
rect 11940 15810 12000 16906
rect 12270 16860 12420 17010
rect 13530 16920 13650 17010
rect 12270 15990 12284 16860
rect 12406 15990 12420 16860
rect 12270 15930 12420 15990
rect 12540 16906 12660 16920
rect 11940 15734 12060 15810
rect 11760 15720 12060 15734
rect 12420 15734 12540 15810
rect 12420 15720 12660 15734
rect 13260 16906 13380 16920
rect 13500 16860 13650 16920
rect 13500 15990 13514 16860
rect 13636 15990 13650 16860
rect 13500 15930 13650 15990
rect 13920 16906 14160 16920
rect 13380 15734 13470 15810
rect 13260 15720 13470 15734
rect 13920 15734 13980 16906
rect 14100 15810 14160 16906
rect 14430 16860 14580 17010
rect 15210 16920 15330 17010
rect 14430 15990 14444 16860
rect 14566 15990 14580 16860
rect 14430 15930 14580 15990
rect 14700 16906 14820 16920
rect 14100 15734 14220 15810
rect 13920 15720 14220 15734
rect 14580 15734 14700 15810
rect 14580 15720 14820 15734
rect 14940 16906 15060 16920
rect 15180 16860 15330 16920
rect 15180 15990 15194 16860
rect 15316 15990 15330 16860
rect 15180 15930 15330 15990
rect 15600 16906 15840 16920
rect 15060 15734 15210 15810
rect 14940 15720 15210 15734
rect 15600 15734 15660 16906
rect 15780 15734 15840 16906
rect 16110 16860 16260 17010
rect 16860 16920 16980 17010
rect 16110 15990 16124 16860
rect 16246 15990 16260 16860
rect 16110 15930 16260 15990
rect 16380 16906 16500 16920
rect 15600 15720 15840 15734
rect 16260 15734 16380 15810
rect 16260 15720 16500 15734
rect 16620 16876 16740 16920
rect 17100 16906 17220 16920
rect 16620 15810 16740 15854
rect 16620 15734 17100 15810
rect 16620 15720 17220 15734
rect 17340 16906 17460 16920
rect 17340 15720 17460 15734
rect 17580 16890 17700 16920
rect 17820 16890 17940 17010
rect 18150 16906 18270 17010
rect 18150 16320 18270 16334
rect 18390 16906 18510 16920
rect 8490 15510 8580 15720
rect 8460 15390 8580 15510
rect 10170 15510 10260 15720
rect 11340 15630 11430 15720
rect 11340 15540 11730 15630
rect 11970 15510 12060 15720
rect 13500 15630 13590 15720
rect 13500 15540 13890 15630
rect 14130 15510 14220 15720
rect 10140 15390 10260 15510
rect 7980 15150 8280 15240
rect 8490 15210 8580 15390
rect 7980 15120 8070 15150
rect 8490 15120 8640 15210
rect 6300 14866 6420 14880
rect 7740 14880 8010 14970
rect 6660 14866 6810 14880
rect 6660 14790 6690 14866
rect 6300 14190 6420 14294
rect 6690 14280 6810 14294
rect 7740 14866 7860 14880
rect 8550 14820 8640 15120
rect 9660 15150 9960 15240
rect 10170 15210 10260 15390
rect 11970 15420 12180 15510
rect 11520 15330 11790 15420
rect 11700 15240 11790 15330
rect 11910 15390 12180 15420
rect 11910 15330 12060 15390
rect 14130 15420 14340 15510
rect 13680 15330 13950 15420
rect 9660 15120 9750 15150
rect 10170 15120 10320 15210
rect 8760 15030 8850 15090
rect 9060 14880 9300 14970
rect 7740 14280 7860 14294
rect 7980 14746 8130 14790
rect 7980 14324 7994 14746
rect 8116 14324 8130 14746
rect 7980 14280 8130 14324
rect 8400 14760 8640 14820
rect 9180 14866 9300 14880
rect 8400 14340 8460 14760
rect 8580 14340 8640 14760
rect 8400 14280 8640 14340
rect 8910 14746 9060 14790
rect 8910 14324 8924 14746
rect 9046 14324 9060 14746
rect 8010 14190 8130 14280
rect 8910 14190 9060 14324
rect 9180 14280 9300 14294
rect 9420 14880 9690 14970
rect 9420 14866 9540 14880
rect 10230 14820 10320 15120
rect 10860 15090 10980 15210
rect 11100 15090 11220 15210
rect 11340 15090 11610 15180
rect 10440 15030 10530 15090
rect 11520 15030 11610 15090
rect 10740 14880 10980 14970
rect 9420 14280 9540 14294
rect 9660 14746 9810 14790
rect 9660 14324 9674 14746
rect 9796 14324 9810 14746
rect 9660 14280 9810 14324
rect 10080 14760 10320 14820
rect 10860 14866 10980 14880
rect 10080 14340 10140 14760
rect 10260 14340 10320 14760
rect 10080 14280 10320 14340
rect 10590 14746 10740 14790
rect 10590 14324 10604 14746
rect 10726 14324 10740 14746
rect 9690 14190 9810 14280
rect 10590 14190 10740 14324
rect 10860 14280 10980 14294
rect 11100 14880 11310 14970
rect 11520 14940 11580 15030
rect 11100 14866 11220 14880
rect 11910 14820 12000 15330
rect 13860 15240 13950 15330
rect 14070 15390 14340 15420
rect 15690 15510 15780 15720
rect 15660 15390 15780 15510
rect 16620 15495 16740 15510
rect 14070 15330 14220 15390
rect 12540 15195 12660 15210
rect 12540 15105 13020 15195
rect 12540 15090 12660 15105
rect 13260 15090 13380 15210
rect 13500 15090 13770 15180
rect 12120 15030 12210 15090
rect 13680 15030 13770 15090
rect 12420 14880 12660 14970
rect 11100 14280 11220 14294
rect 11340 14746 11490 14790
rect 11340 14324 11354 14746
rect 11476 14324 11490 14746
rect 11340 14280 11490 14324
rect 11760 14760 12000 14820
rect 12540 14866 12660 14880
rect 11760 14340 11820 14760
rect 11940 14340 12000 14760
rect 11760 14280 12000 14340
rect 12270 14746 12420 14790
rect 12270 14324 12284 14746
rect 12406 14324 12420 14746
rect 11370 14190 11490 14280
rect 12270 14190 12420 14324
rect 12540 14280 12660 14294
rect 13260 14880 13470 14970
rect 13680 14940 13740 15030
rect 13260 14866 13380 14880
rect 14070 14820 14160 15330
rect 15180 15150 15480 15240
rect 15690 15210 15780 15390
rect 16395 15450 16740 15495
rect 17340 15510 17430 15720
rect 16395 15420 16860 15450
rect 17100 15420 17460 15510
rect 16395 15405 16740 15420
rect 16395 15210 16485 15405
rect 16620 15390 16740 15405
rect 15180 15120 15270 15150
rect 15690 15120 15840 15210
rect 14280 15030 14370 15090
rect 14580 14880 14820 14970
rect 13260 14280 13380 14294
rect 13500 14746 13650 14790
rect 13500 14324 13514 14746
rect 13636 14324 13650 14746
rect 13500 14280 13650 14324
rect 13920 14760 14160 14820
rect 14700 14866 14820 14880
rect 13920 14340 13980 14760
rect 14100 14340 14160 14760
rect 13920 14280 14160 14340
rect 14430 14746 14580 14790
rect 14430 14324 14444 14746
rect 14566 14324 14580 14746
rect 13530 14190 13650 14280
rect 14430 14190 14580 14324
rect 14700 14280 14820 14294
rect 14940 14880 15210 14970
rect 14940 14866 15060 14880
rect 15750 14820 15840 15120
rect 16380 15195 16500 15210
rect 16620 15195 16740 15210
rect 16380 15105 16740 15195
rect 16380 15090 16500 15105
rect 16620 15090 16740 15105
rect 15960 15030 16050 15090
rect 16260 14880 16500 14970
rect 17100 14880 17190 15420
rect 17340 15390 17460 15420
rect 17340 14895 17460 14910
rect 17580 14895 17700 16320
rect 18180 15810 18270 15990
rect 18060 15795 18270 15810
rect 17940 15720 18270 15795
rect 18360 15734 18390 15810
rect 18360 15720 18510 15734
rect 18780 16906 18900 17010
rect 19260 16906 19380 17010
rect 19260 16320 19380 16334
rect 19500 16906 19620 16920
rect 18780 15720 18900 15734
rect 17940 15705 18180 15720
rect 18060 15690 18180 15705
rect 18360 15210 18450 15720
rect 18060 15090 18450 15210
rect 18780 15180 18900 15210
rect 18660 15150 18900 15180
rect 14940 14280 15060 14294
rect 15180 14746 15330 14790
rect 15180 14324 15194 14746
rect 15316 14324 15330 14746
rect 15180 14280 15330 14324
rect 15600 14760 15840 14820
rect 16380 14866 16500 14880
rect 15600 14340 15660 14760
rect 15780 14340 15840 14760
rect 15600 14280 15840 14340
rect 16110 14746 16260 14790
rect 16110 14324 16124 14746
rect 16246 14324 16260 14746
rect 15210 14190 15330 14280
rect 16110 14190 16260 14324
rect 16380 14280 16500 14294
rect 16710 14866 16830 14880
rect 16710 14190 16830 14294
rect 17100 14866 17220 14880
rect 17340 14805 17700 14895
rect 17340 14790 17460 14805
rect 17100 14280 17220 14294
rect 17340 14566 17460 14580
rect 17340 14190 17460 14294
rect 17580 14550 17700 14805
rect 17820 14895 17940 14910
rect 18075 14895 18180 15090
rect 18780 15090 18900 15150
rect 17820 14866 18180 14895
rect 18330 14880 18870 14940
rect 19500 14910 19620 16334
rect 19740 16906 19860 17010
rect 19740 16320 19860 16334
rect 20700 16906 20820 17010
rect 19740 15795 19860 15810
rect 19740 15705 20460 15795
rect 19740 15690 19860 15705
rect 20700 15720 20820 15734
rect 21090 16906 21210 16920
rect 21330 16906 21450 17010
rect 21330 16320 21450 16334
rect 22230 16906 22350 17010
rect 22230 16320 22350 16334
rect 22470 16906 22590 16920
rect 21330 15810 21420 15990
rect 22260 15810 22350 15990
rect 21210 15734 21240 15810
rect 21090 15720 21240 15734
rect 21330 15795 21540 15810
rect 21330 15720 21660 15795
rect 20940 15495 21060 15510
rect 20100 15405 21060 15495
rect 20940 15390 21060 15405
rect 21150 15210 21240 15720
rect 21420 15705 21660 15720
rect 21420 15690 21540 15705
rect 22140 15720 22350 15810
rect 22440 15734 22470 15810
rect 22440 15720 22590 15734
rect 22860 16906 22980 17010
rect 23580 16906 23700 17010
rect 23580 16320 23700 16334
rect 23820 16906 23940 16920
rect 22860 15720 22980 15734
rect 22140 15690 22260 15720
rect 22440 15210 22530 15720
rect 22620 15390 22740 15510
rect 23820 15495 23940 16334
rect 24060 16906 24180 17010
rect 24060 16320 24180 16334
rect 24780 16906 24900 17010
rect 24780 16320 24900 16334
rect 25020 16906 25140 16920
rect 24780 15795 24900 15810
rect 24315 15705 24900 15795
rect 24315 15495 24405 15705
rect 24780 15690 24900 15705
rect 23820 15405 24405 15495
rect 21150 15195 21540 15210
rect 20820 15150 20940 15180
rect 21150 15105 21900 15195
rect 21150 15090 21540 15105
rect 22140 15090 22530 15210
rect 22860 15195 22980 15210
rect 23580 15195 23700 15210
rect 22860 15180 23700 15195
rect 22740 15150 23700 15180
rect 17820 14805 18060 14866
rect 17820 14790 17940 14805
rect 17820 14550 17940 14580
rect 18060 14280 18180 14294
rect 18300 14866 18900 14880
rect 18420 14850 18780 14866
rect 18300 14280 18420 14294
rect 18540 14730 18660 14760
rect 17820 14190 17940 14280
rect 18540 14190 18660 14310
rect 18780 14280 18900 14294
rect 19260 14866 19380 14880
rect 20730 14880 21270 14940
rect 21420 14880 21510 15090
rect 22170 14880 22260 15090
rect 22860 15105 23700 15150
rect 22860 15090 22980 15105
rect 23580 15090 23700 15105
rect 22410 14880 22950 14940
rect 23820 14880 23940 15405
rect 25020 14880 25140 16334
rect 25260 16906 25380 17010
rect 25260 16320 25380 16334
rect 25740 16906 25860 16920
rect 25980 16860 26130 17010
rect 26910 16920 27030 17010
rect 25980 15990 25994 16860
rect 26116 15990 26130 16860
rect 25980 15930 26130 15990
rect 26400 16906 26640 16920
rect 25860 15734 25980 15810
rect 25740 15720 25980 15734
rect 26400 15734 26460 16906
rect 26580 15734 26640 16906
rect 26910 16860 27060 16920
rect 26910 15990 26924 16860
rect 27046 15990 27060 16860
rect 26910 15930 27060 15990
rect 27180 16906 27300 16920
rect 26400 15720 26640 15734
rect 27030 15734 27180 15810
rect 27900 16906 28020 17010
rect 27900 16320 28020 16334
rect 28140 16906 28260 16920
rect 27030 15720 27300 15734
rect 26460 15510 26550 15720
rect 26460 15390 26580 15510
rect 28140 15495 28260 16334
rect 28380 16906 28500 17010
rect 28380 16320 28500 16334
rect 29100 16906 29220 17010
rect 29100 16320 29220 16334
rect 29340 16906 29460 16920
rect 27675 15405 28260 15495
rect 26460 15210 26550 15390
rect 25740 15195 25860 15210
rect 25620 15105 25860 15195
rect 25740 15090 25860 15105
rect 26190 15030 26280 15090
rect 26400 15120 26550 15210
rect 26760 15150 27060 15240
rect 26970 15120 27060 15150
rect 25740 14880 25980 14970
rect 19620 14866 19770 14880
rect 19620 14790 19650 14866
rect 19260 14190 19380 14294
rect 19650 14280 19770 14294
rect 20700 14866 21300 14880
rect 20820 14850 21180 14866
rect 20700 14280 20820 14294
rect 20940 14730 21060 14760
rect 20940 14190 21060 14310
rect 21180 14280 21300 14294
rect 21420 14866 21540 14880
rect 22140 14866 22260 14880
rect 22020 14505 22140 14595
rect 21420 14280 21540 14294
rect 22140 14280 22260 14294
rect 22380 14866 22980 14880
rect 22500 14850 22860 14866
rect 22380 14280 22500 14294
rect 22620 14730 22740 14760
rect 22620 14190 22740 14310
rect 22860 14280 22980 14294
rect 23580 14866 23700 14880
rect 23820 14866 24090 14880
rect 23820 14790 23970 14866
rect 23580 14190 23700 14294
rect 23970 14280 24090 14294
rect 24870 14866 25140 14880
rect 24990 14790 25140 14866
rect 25260 14866 25380 14880
rect 24870 14280 24990 14294
rect 25260 14190 25380 14294
rect 25740 14866 25860 14880
rect 26400 14820 26490 15120
rect 27180 15195 27300 15210
rect 27675 15195 27765 15405
rect 27180 15105 27765 15195
rect 27180 15090 27300 15105
rect 27030 14880 27300 14970
rect 28140 14880 28260 15405
rect 29340 15495 29460 16334
rect 29580 16906 29700 17010
rect 29580 16320 29700 16334
rect 30300 16906 30420 16920
rect 29580 15795 29700 15810
rect 30060 15795 30180 15810
rect 29580 15705 30180 15795
rect 30540 16860 30690 17010
rect 31470 16920 31590 17010
rect 30540 15990 30554 16860
rect 30676 15990 30690 16860
rect 30540 15930 30690 15990
rect 30960 16906 31200 16920
rect 30420 15734 30540 15810
rect 30300 15720 30540 15734
rect 30960 15734 31020 16906
rect 31140 15734 31200 16906
rect 31470 16860 31620 16920
rect 31470 15990 31484 16860
rect 31606 15990 31620 16860
rect 31470 15930 31620 15990
rect 31740 16906 31860 16920
rect 30960 15720 31200 15734
rect 31590 15734 31740 15810
rect 32220 16906 32340 17010
rect 32220 16320 32340 16334
rect 32460 16906 32580 16920
rect 31590 15720 31860 15734
rect 31980 15795 32100 15810
rect 32220 15795 32340 15810
rect 29580 15690 29700 15705
rect 30060 15690 30180 15705
rect 28740 15405 29460 15495
rect 28500 15105 29100 15195
rect 29340 14880 29460 15405
rect 31020 15510 31110 15720
rect 31980 15705 32340 15795
rect 31980 15690 32100 15705
rect 32220 15690 32340 15705
rect 31020 15390 31140 15510
rect 31020 15210 31110 15390
rect 30750 15030 30840 15090
rect 30960 15120 31110 15210
rect 31320 15150 31620 15240
rect 31530 15120 31620 15150
rect 30300 14880 30540 14970
rect 27180 14866 27300 14880
rect 25740 14280 25860 14294
rect 25980 14746 26130 14790
rect 25980 14324 25994 14746
rect 26116 14324 26130 14746
rect 25980 14190 26130 14324
rect 26400 14760 26640 14820
rect 26400 14340 26460 14760
rect 26580 14340 26640 14760
rect 26400 14280 26640 14340
rect 26910 14746 27060 14790
rect 26910 14324 26924 14746
rect 27046 14324 27060 14746
rect 26910 14280 27060 14324
rect 27180 14280 27300 14294
rect 27900 14866 28020 14880
rect 28140 14866 28410 14880
rect 28140 14790 28290 14866
rect 26910 14190 27030 14280
rect 27900 14190 28020 14294
rect 28290 14280 28410 14294
rect 29100 14866 29220 14880
rect 29340 14866 29610 14880
rect 29340 14790 29490 14866
rect 29100 14190 29220 14294
rect 29490 14280 29610 14294
rect 30300 14866 30420 14880
rect 30960 14820 31050 15120
rect 31590 14880 31860 14970
rect 32460 14880 32580 16334
rect 32700 16906 32820 17010
rect 32700 16320 32820 16334
rect 33180 16906 33300 17010
rect 33180 16320 33300 16334
rect 33420 16906 33540 16920
rect 32700 15195 32820 15210
rect 32700 15105 32940 15195
rect 32700 15090 32820 15105
rect 33420 14895 33540 16334
rect 33660 16906 33780 17010
rect 33660 16320 33780 16334
rect 34620 16906 34740 17010
rect 34620 16320 34740 16334
rect 34860 16906 34980 16920
rect 33780 15105 34620 15195
rect 31740 14866 31860 14880
rect 30300 14280 30420 14294
rect 30540 14746 30690 14790
rect 30540 14324 30554 14746
rect 30676 14324 30690 14746
rect 30540 14190 30690 14324
rect 30960 14760 31200 14820
rect 30960 14340 31020 14760
rect 31140 14340 31200 14760
rect 30960 14280 31200 14340
rect 31470 14746 31620 14790
rect 31470 14324 31484 14746
rect 31606 14324 31620 14746
rect 31470 14280 31620 14324
rect 31740 14280 31860 14294
rect 32310 14866 32580 14880
rect 32430 14790 32580 14866
rect 32700 14866 32820 14880
rect 32310 14280 32430 14294
rect 31470 14190 31590 14280
rect 32700 14190 32820 14294
rect 33180 14866 33300 14880
rect 33420 14866 34380 14895
rect 33420 14790 33570 14866
rect 33180 14190 33300 14294
rect 33690 14805 34380 14866
rect 34860 14895 34980 16334
rect 35100 16906 35220 17010
rect 35100 16320 35220 16334
rect 36060 16906 36180 17010
rect 35100 15795 35220 15810
rect 35100 15705 35580 15795
rect 35100 15690 35220 15705
rect 35820 15795 35940 15810
rect 35700 15705 35940 15795
rect 36060 15720 36180 15734
rect 36450 16906 36570 16920
rect 36690 16906 36810 17010
rect 36690 16320 36810 16334
rect 37740 16906 37860 17010
rect 37740 16320 37860 16334
rect 37980 16906 38100 16920
rect 36690 15810 36780 15990
rect 36570 15734 36600 15810
rect 36450 15720 36600 15734
rect 36690 15795 36900 15810
rect 36690 15720 37740 15795
rect 35820 15690 35940 15705
rect 36300 15390 36420 15510
rect 36510 15210 36600 15720
rect 36780 15705 37740 15720
rect 36780 15690 36900 15705
rect 35100 15195 35220 15210
rect 36060 15195 36180 15210
rect 35100 15180 36180 15195
rect 35100 15150 36300 15180
rect 35100 15105 36180 15150
rect 35100 15090 35220 15105
rect 36060 15090 36180 15105
rect 36510 15090 36900 15210
rect 37020 15195 37140 15210
rect 37020 15105 37740 15195
rect 37020 15090 37140 15105
rect 34620 14866 34740 14880
rect 33570 14280 33690 14294
rect 34860 14866 35820 14895
rect 34860 14790 35010 14866
rect 34620 14190 34740 14294
rect 35130 14805 35820 14866
rect 36090 14880 36630 14940
rect 36780 14880 36870 15090
rect 37980 14880 38100 16334
rect 38220 16906 38340 17010
rect 38220 16320 38340 16334
rect 38700 16906 38820 16920
rect 38940 16860 39090 17010
rect 39870 16920 39990 17010
rect 41850 16920 41970 17010
rect 38940 15990 38954 16860
rect 39076 15990 39090 16860
rect 38940 15930 39090 15990
rect 39360 16906 39600 16920
rect 38820 15734 38940 15810
rect 38700 15720 38940 15734
rect 39360 15734 39420 16906
rect 39540 15734 39600 16906
rect 39870 16860 40020 16920
rect 39870 15990 39884 16860
rect 40006 15990 40020 16860
rect 39870 15930 40020 15990
rect 40140 16906 40260 16920
rect 39360 15720 39600 15734
rect 39990 15734 40140 15810
rect 39990 15720 40260 15734
rect 41580 16906 41700 16920
rect 41820 16860 41970 16920
rect 41820 15990 41834 16860
rect 41956 15990 41970 16860
rect 41820 15930 41970 15990
rect 42240 16906 42480 16920
rect 41700 15734 41850 15810
rect 41580 15720 41850 15734
rect 42240 15734 42300 16906
rect 42420 15734 42480 16906
rect 42750 16860 42900 17010
rect 42750 15990 42764 16860
rect 42886 15990 42900 16860
rect 42750 15930 42900 15990
rect 43020 16906 43140 16920
rect 42240 15720 42480 15734
rect 42900 15734 43020 15810
rect 42900 15720 43140 15734
rect 44460 16906 44580 17010
rect 44460 15720 44580 15734
rect 44850 16906 44970 16920
rect 45090 16906 45210 17010
rect 45090 16320 45210 16334
rect 46140 16906 46260 17010
rect 46140 16320 46260 16334
rect 46380 16906 46500 16920
rect 45090 15810 45180 15990
rect 44970 15734 45000 15810
rect 44850 15720 45000 15734
rect 45090 15795 45300 15810
rect 46380 15795 46500 16334
rect 46620 16906 46740 17010
rect 46620 16320 46740 16334
rect 47580 16906 47700 17010
rect 47580 16320 47700 16334
rect 47820 16906 47940 16920
rect 45090 15720 46500 15795
rect 39420 15510 39510 15720
rect 39420 15495 39540 15510
rect 38820 15405 39540 15495
rect 39420 15390 39540 15405
rect 42330 15510 42420 15720
rect 42300 15390 42420 15510
rect 39420 15210 39510 15390
rect 38700 15195 38820 15210
rect 38580 15105 38820 15195
rect 38700 15090 38820 15105
rect 39150 15030 39240 15090
rect 39360 15120 39510 15210
rect 39720 15150 40020 15240
rect 39930 15120 40020 15150
rect 38700 14880 38940 14970
rect 36060 14866 36660 14880
rect 35010 14280 35130 14294
rect 36180 14850 36540 14866
rect 36060 14280 36180 14294
rect 36300 14730 36420 14760
rect 36300 14190 36420 14310
rect 36540 14280 36660 14294
rect 36780 14866 36900 14880
rect 36780 14280 36900 14294
rect 37740 14866 37860 14880
rect 37980 14866 38250 14880
rect 37980 14790 38130 14866
rect 37740 14190 37860 14294
rect 38130 14280 38250 14294
rect 38700 14866 38820 14880
rect 39360 14820 39450 15120
rect 40140 15195 40260 15210
rect 40140 15105 41340 15195
rect 40140 15090 40260 15105
rect 41820 15150 42120 15240
rect 42330 15210 42420 15390
rect 44910 15210 45000 15720
rect 45180 15705 46500 15720
rect 45180 15690 45300 15705
rect 41820 15120 41910 15150
rect 42330 15120 42480 15210
rect 39990 14880 40260 14970
rect 40140 14866 40260 14880
rect 38700 14280 38820 14294
rect 38940 14746 39090 14790
rect 38940 14324 38954 14746
rect 39076 14324 39090 14746
rect 38940 14190 39090 14324
rect 39360 14760 39600 14820
rect 39360 14340 39420 14760
rect 39540 14340 39600 14760
rect 39360 14280 39600 14340
rect 39870 14746 40020 14790
rect 39870 14324 39884 14746
rect 40006 14324 40020 14746
rect 39870 14280 40020 14324
rect 40140 14280 40260 14294
rect 41580 14880 41850 14970
rect 41580 14866 41700 14880
rect 42390 14820 42480 15120
rect 43020 15090 43140 15210
rect 43620 15105 44460 15195
rect 44580 15150 44700 15180
rect 42600 15030 42690 15090
rect 44910 15090 45180 15210
rect 45420 15195 45540 15210
rect 46140 15195 46260 15210
rect 45420 15105 46260 15195
rect 45420 15090 45540 15105
rect 46140 15090 46260 15105
rect 42900 14880 43140 14970
rect 44490 14880 45030 14940
rect 45180 14880 45270 15090
rect 46380 14880 46500 15705
rect 46620 15690 46740 15810
rect 47580 15795 47700 15810
rect 46980 15705 47700 15795
rect 47580 15690 47700 15705
rect 47820 14880 47940 16334
rect 48060 16906 48180 17010
rect 48060 16320 48180 16334
rect 49020 16906 49140 17010
rect 49020 15720 49140 15734
rect 49410 16906 49530 16920
rect 49650 16906 49770 17010
rect 49650 16320 49770 16334
rect 49650 15810 49740 15990
rect 49530 15734 49560 15810
rect 49410 15720 49560 15734
rect 49650 15795 49860 15810
rect 49650 15720 49980 15795
rect 49260 15390 49380 15510
rect 49470 15210 49560 15720
rect 49740 15705 49980 15720
rect 49740 15690 49860 15705
rect 49020 15195 49140 15210
rect 48900 15180 49140 15195
rect 48900 15150 49260 15180
rect 48900 15105 49140 15150
rect 49020 15090 49140 15105
rect 49470 15090 49860 15210
rect 49050 14880 49590 14940
rect 49740 14880 49830 15090
rect 41580 14280 41700 14294
rect 41820 14746 41970 14790
rect 41820 14324 41834 14746
rect 41956 14324 41970 14746
rect 41820 14280 41970 14324
rect 42240 14760 42480 14820
rect 43020 14866 43140 14880
rect 42240 14340 42300 14760
rect 42420 14340 42480 14760
rect 42240 14280 42480 14340
rect 42750 14746 42900 14790
rect 42750 14324 42764 14746
rect 42886 14324 42900 14746
rect 39870 14190 39990 14280
rect 41850 14190 41970 14280
rect 42750 14190 42900 14324
rect 43020 14280 43140 14294
rect 44460 14866 45060 14880
rect 44580 14850 44940 14866
rect 44460 14280 44580 14294
rect 44700 14730 44820 14760
rect 44700 14190 44820 14310
rect 44940 14280 45060 14294
rect 45180 14866 45300 14880
rect 45180 14280 45300 14294
rect 46140 14866 46260 14880
rect 46380 14866 46650 14880
rect 46380 14790 46530 14866
rect 46140 14190 46260 14294
rect 46530 14280 46650 14294
rect 47670 14866 47940 14880
rect 47790 14790 47940 14866
rect 48060 14866 48180 14880
rect 47670 14280 47790 14294
rect 48060 14190 48180 14294
rect 49020 14866 49620 14880
rect 49140 14850 49500 14866
rect 49020 14280 49140 14294
rect 49260 14730 49380 14760
rect 49260 14190 49380 14310
rect 49500 14280 49620 14294
rect 49740 14866 49860 14880
rect 49740 14280 49860 14294
rect 3135 14160 52260 14190
rect 3135 14040 3194 14160
rect 4066 14040 5220 14160
rect 5340 14040 5460 14160
rect 5580 14040 5700 14160
rect 5820 14040 5940 14160
rect 6060 14040 6180 14160
rect 6300 14040 6420 14160
rect 6540 14040 6660 14160
rect 6780 14040 6900 14160
rect 7020 14040 7140 14160
rect 7260 14040 7380 14160
rect 7500 14040 7620 14160
rect 7740 14040 7860 14160
rect 7980 14040 8100 14160
rect 8220 14040 8340 14160
rect 8460 14040 8580 14160
rect 8700 14040 8820 14160
rect 8940 14040 9060 14160
rect 9180 14040 9300 14160
rect 9420 14040 9780 14160
rect 9900 14040 10020 14160
rect 10140 14040 10260 14160
rect 10380 14040 10500 14160
rect 10620 14040 10740 14160
rect 10860 14040 10980 14160
rect 11100 14040 11220 14160
rect 11340 14040 11460 14160
rect 11580 14040 11700 14160
rect 11820 14040 11940 14160
rect 12060 14040 12420 14160
rect 12540 14040 12660 14160
rect 12780 14040 12900 14160
rect 13020 14040 13140 14160
rect 13260 14040 13380 14160
rect 13500 14040 13620 14160
rect 13740 14040 13860 14160
rect 13980 14040 14100 14160
rect 14220 14040 14340 14160
rect 14460 14040 14580 14160
rect 14700 14040 14820 14160
rect 14940 14040 15060 14160
rect 15180 14040 15300 14160
rect 15420 14040 15540 14160
rect 15660 14040 15780 14160
rect 15900 14040 16260 14160
rect 16380 14040 16500 14160
rect 16620 14040 16980 14160
rect 17100 14040 17460 14160
rect 17580 14040 17940 14160
rect 18060 14040 18420 14160
rect 18540 14040 18900 14160
rect 19020 14040 19140 14160
rect 19260 14040 19380 14160
rect 19500 14040 19620 14160
rect 19740 14040 19860 14160
rect 19980 14040 20100 14160
rect 20220 14040 20340 14160
rect 20460 14040 20580 14160
rect 20700 14040 20820 14160
rect 20940 14040 21060 14160
rect 21180 14040 21300 14160
rect 21420 14040 21540 14160
rect 21660 14040 21780 14160
rect 21900 14040 22020 14160
rect 22140 14040 22260 14160
rect 22380 14040 22500 14160
rect 22620 14040 22740 14160
rect 22860 14040 22980 14160
rect 23100 14040 23220 14160
rect 23340 14040 23460 14160
rect 23580 14040 23700 14160
rect 23820 14040 23940 14160
rect 24060 14040 24180 14160
rect 24300 14040 24420 14160
rect 24540 14040 24660 14160
rect 24780 14040 24900 14160
rect 25020 14040 25380 14160
rect 25500 14040 25620 14160
rect 25740 14040 25860 14160
rect 25980 14040 26100 14160
rect 26220 14040 26340 14160
rect 26460 14040 26580 14160
rect 26700 14040 26820 14160
rect 26940 14040 27060 14160
rect 27180 14040 27300 14160
rect 27420 14040 27540 14160
rect 27660 14040 27780 14160
rect 27900 14040 28020 14160
rect 28140 14040 28260 14160
rect 28380 14040 28500 14160
rect 28620 14040 28740 14160
rect 28860 14040 28980 14160
rect 29100 14040 29460 14160
rect 29580 14040 29700 14160
rect 29820 14040 29940 14160
rect 30060 14040 30180 14160
rect 30300 14040 30420 14160
rect 30540 14040 30660 14160
rect 30780 14040 30900 14160
rect 31020 14040 31140 14160
rect 31260 14040 31380 14160
rect 31500 14040 31620 14160
rect 31740 14040 31860 14160
rect 31980 14040 32100 14160
rect 32220 14040 32340 14160
rect 32460 14040 32580 14160
rect 32700 14040 32820 14160
rect 32940 14040 33060 14160
rect 33180 14040 33300 14160
rect 33420 14040 33540 14160
rect 33660 14040 33780 14160
rect 33900 14040 34020 14160
rect 34140 14040 34260 14160
rect 34380 14040 34500 14160
rect 34620 14040 34980 14160
rect 35100 14040 35220 14160
rect 35340 14040 35460 14160
rect 35580 14040 35700 14160
rect 35820 14040 35940 14160
rect 36060 14040 36420 14160
rect 36540 14040 36660 14160
rect 36780 14040 36900 14160
rect 37020 14040 37140 14160
rect 37260 14040 37380 14160
rect 37500 14040 37620 14160
rect 37740 14040 37860 14160
rect 37980 14040 38100 14160
rect 38220 14040 38340 14160
rect 38460 14040 38580 14160
rect 38700 14040 38820 14160
rect 38940 14040 39300 14160
rect 39420 14040 39540 14160
rect 39660 14040 39780 14160
rect 39900 14040 40020 14160
rect 40140 14040 40260 14160
rect 40380 14040 40500 14160
rect 40620 14040 40740 14160
rect 40860 14040 40980 14160
rect 41100 14040 41220 14160
rect 41340 14040 41460 14160
rect 41580 14040 41940 14160
rect 42060 14040 42420 14160
rect 42540 14040 42660 14160
rect 42780 14040 42900 14160
rect 43020 14040 43140 14160
rect 43260 14040 43380 14160
rect 43500 14040 43620 14160
rect 43740 14040 43860 14160
rect 43980 14040 44100 14160
rect 44220 14040 44340 14160
rect 44460 14040 44820 14160
rect 44940 14040 45300 14160
rect 45420 14040 45540 14160
rect 45660 14040 45780 14160
rect 45900 14040 46020 14160
rect 46140 14040 46500 14160
rect 46620 14040 46740 14160
rect 46860 14040 46980 14160
rect 47100 14040 47220 14160
rect 47340 14040 47460 14160
rect 47580 14040 47700 14160
rect 47820 14040 47940 14160
rect 48060 14040 48180 14160
rect 48300 14040 48420 14160
rect 48540 14040 48660 14160
rect 48780 14040 48900 14160
rect 49020 14040 49140 14160
rect 49260 14040 49380 14160
rect 49500 14040 49860 14160
rect 49980 14040 50100 14160
rect 50220 14040 51330 14160
rect 52200 14040 52260 14160
rect 3135 14010 52260 14040
rect 6870 13906 6990 13920
rect 5700 13334 6870 13395
rect 7260 13906 7380 14010
rect 6990 13334 7140 13410
rect 5700 13305 7140 13334
rect 7260 13320 7380 13334
rect 8940 13906 9060 13920
rect 9180 13890 9300 14010
rect 9180 13440 9300 13470
rect 9420 13906 10020 13920
rect 9060 13334 9420 13350
rect 9540 13830 9900 13906
rect 8940 13320 9540 13334
rect 9900 13320 10020 13334
rect 10860 13906 10980 14010
rect 11250 13906 11370 13920
rect 10860 13320 10980 13334
rect 11100 13334 11250 13410
rect 12060 13906 12180 13920
rect 11700 13605 12060 13695
rect 11100 13320 11370 13334
rect 12060 13320 12180 13334
rect 12300 13906 12420 13920
rect 12540 13890 12660 14010
rect 12540 13440 12660 13470
rect 12780 13906 12900 13920
rect 12420 13334 12780 13350
rect 12300 13320 12900 13334
rect 15900 13906 16020 14010
rect 16290 13906 16410 13920
rect 15900 13320 16020 13334
rect 16140 13334 16290 13410
rect 16140 13320 16410 13334
rect 16620 13906 16740 13920
rect 16620 13320 16740 13334
rect 16860 13906 16980 13920
rect 17100 13890 17220 14010
rect 17850 13920 17970 14010
rect 17100 13440 17220 13470
rect 17340 13906 17460 13920
rect 16980 13334 17340 13350
rect 16860 13320 17460 13334
rect 17580 13906 17700 13920
rect 17820 13876 17970 13920
rect 17820 13454 17834 13876
rect 17956 13454 17970 13876
rect 17820 13410 17970 13454
rect 18240 13860 18480 13920
rect 18240 13440 18300 13860
rect 18420 13440 18480 13860
rect 18240 13380 18480 13440
rect 18750 13876 18900 14010
rect 18750 13454 18764 13876
rect 18886 13454 18900 13876
rect 18750 13410 18900 13454
rect 19020 13906 19140 13920
rect 17580 13320 17700 13334
rect 6780 12495 6900 12510
rect 6660 12405 6900 12495
rect 6780 12390 6900 12405
rect 6780 11866 6900 11880
rect 6780 11190 6900 11294
rect 7020 11866 7140 13305
rect 8970 13260 9510 13320
rect 7260 13095 7380 13110
rect 7260 13005 7740 13095
rect 7260 12990 7380 13005
rect 8220 13095 8340 13110
rect 7860 13005 8340 13095
rect 8220 12990 8340 13005
rect 8940 13095 9060 13110
rect 8580 13050 9060 13095
rect 9690 13110 9780 13320
rect 8580 13020 9180 13050
rect 9420 13020 9780 13110
rect 8580 13005 9060 13020
rect 8940 12990 9060 13005
rect 9420 12990 9540 13020
rect 10860 12990 10980 13110
rect 9420 12480 9510 12990
rect 8940 12466 9060 12480
rect 7020 11280 7140 11294
rect 7260 11866 7380 11880
rect 7260 11190 7380 11294
rect 8940 11190 9060 11294
rect 9330 12466 9630 12480
rect 9330 11294 9344 12466
rect 9616 11294 9630 12466
rect 9330 11280 9630 11294
rect 9900 12466 10020 12480
rect 9900 11190 10020 11294
rect 10860 11866 10980 11880
rect 10860 11190 10980 11294
rect 11100 11866 11220 13320
rect 12090 13110 12180 13320
rect 12330 13260 12870 13320
rect 12060 12990 12450 13110
rect 12780 13050 12900 13110
rect 12660 13020 12900 13050
rect 12780 12990 12900 13020
rect 11340 12390 11460 12510
rect 12060 12495 12180 12510
rect 11700 12480 12180 12495
rect 12360 12480 12450 12990
rect 16140 12795 16260 13320
rect 16650 13110 16740 13320
rect 16890 13260 17430 13320
rect 17580 13230 17850 13320
rect 16620 12990 17010 13110
rect 17220 13020 17340 13050
rect 17580 13095 17700 13110
rect 17460 13005 17700 13095
rect 17580 12990 17700 13005
rect 18390 13080 18480 13380
rect 19020 13320 19140 13334
rect 18900 13230 19140 13320
rect 19260 13906 19380 13920
rect 19500 13876 19650 14010
rect 20430 13920 20550 14010
rect 22170 13920 22290 14010
rect 19500 13454 19514 13876
rect 19636 13454 19650 13876
rect 19500 13410 19650 13454
rect 19920 13860 20160 13920
rect 19920 13440 19980 13860
rect 20100 13440 20160 13860
rect 19260 13320 19380 13334
rect 19920 13380 20160 13440
rect 20430 13876 20580 13920
rect 20430 13454 20444 13876
rect 20566 13454 20580 13876
rect 20430 13410 20580 13454
rect 20700 13906 20820 13920
rect 19260 13230 19500 13320
rect 17820 13050 17910 13080
rect 16140 12705 16725 12795
rect 11700 12405 12270 12480
rect 12060 12390 12270 12405
rect 12360 12466 12510 12480
rect 12360 12390 12390 12466
rect 12180 12210 12270 12390
rect 11100 11280 11220 11294
rect 11340 11866 11460 11880
rect 11340 11190 11460 11294
rect 12150 11866 12270 11880
rect 12150 11190 12270 11294
rect 12390 11280 12510 11294
rect 12780 12466 12900 12480
rect 12780 11190 12900 11294
rect 15900 11866 16020 11880
rect 15900 11190 16020 11294
rect 16140 11866 16260 12705
rect 16635 12510 16725 12705
rect 16620 12480 16740 12510
rect 16920 12480 17010 12990
rect 17820 12960 18120 13050
rect 18330 12990 18480 13080
rect 18600 13110 18690 13170
rect 19710 13110 19800 13170
rect 19020 12990 19140 13110
rect 19260 12990 19380 13110
rect 18330 12810 18420 12990
rect 18300 12795 18420 12810
rect 19275 12795 19365 12990
rect 19920 12870 20010 13380
rect 20700 13320 20820 13334
rect 20340 13170 20400 13260
rect 20610 13230 20820 13320
rect 21900 13906 22020 13920
rect 22140 13876 22290 13920
rect 22140 13454 22154 13876
rect 22276 13454 22290 13876
rect 22140 13410 22290 13454
rect 22560 13860 22800 13920
rect 22560 13440 22620 13860
rect 22740 13440 22800 13860
rect 22560 13380 22800 13440
rect 23070 13876 23220 14010
rect 23070 13454 23084 13876
rect 23206 13454 23220 13876
rect 23070 13410 23220 13454
rect 23340 13906 23460 13920
rect 21900 13320 22020 13334
rect 21900 13230 22110 13320
rect 20310 13110 20400 13170
rect 22320 13170 22380 13260
rect 22320 13110 22410 13170
rect 20310 13020 20580 13110
rect 20700 12990 20820 13110
rect 21900 12990 22020 13110
rect 22140 13020 22410 13110
rect 19860 12810 20010 12870
rect 18300 12705 19365 12795
rect 19740 12780 20010 12810
rect 20130 12870 20220 12960
rect 22500 12870 22590 12960
rect 20130 12780 20400 12870
rect 18300 12690 18420 12705
rect 19740 12690 19950 12780
rect 22320 12780 22590 12870
rect 22710 12870 22800 13380
rect 23340 13320 23460 13334
rect 25020 13906 25140 13920
rect 25260 13890 25380 14010
rect 25260 13440 25380 13470
rect 25500 13906 25620 13920
rect 25140 13334 25500 13350
rect 25020 13320 25620 13334
rect 25740 13906 25860 13920
rect 25740 13320 25860 13334
rect 26700 13906 26820 14010
rect 27090 13906 27210 13920
rect 26700 13320 26820 13334
rect 26940 13334 27090 13410
rect 26940 13320 27210 13334
rect 29100 13906 29220 13920
rect 29340 13890 29460 14010
rect 29340 13440 29460 13470
rect 29580 13906 29700 13920
rect 29220 13334 29580 13350
rect 29100 13320 29700 13334
rect 29820 13906 29940 13920
rect 29820 13320 29940 13334
rect 30300 13906 30420 13920
rect 30300 13320 30420 13334
rect 30540 13906 30660 13920
rect 30780 13890 30900 14010
rect 30780 13440 30900 13470
rect 31020 13906 31140 13920
rect 30660 13334 31020 13350
rect 30540 13320 31140 13334
rect 32070 13906 32190 13920
rect 32460 13906 32580 14010
rect 33210 13920 33330 14010
rect 32190 13334 32340 13410
rect 32070 13320 32340 13334
rect 32460 13320 32580 13334
rect 32940 13906 33060 13920
rect 33180 13876 33330 13920
rect 33180 13454 33194 13876
rect 33316 13454 33330 13876
rect 33180 13410 33330 13454
rect 33600 13860 33840 13920
rect 33600 13440 33660 13860
rect 33780 13440 33840 13860
rect 33600 13380 33840 13440
rect 34110 13876 34260 14010
rect 34110 13454 34124 13876
rect 34246 13454 34260 13876
rect 34110 13410 34260 13454
rect 34380 13906 34500 13920
rect 32940 13320 33060 13334
rect 23220 13230 23460 13320
rect 25050 13260 25590 13320
rect 22920 13110 23010 13170
rect 23340 13095 23460 13110
rect 24780 13095 24900 13110
rect 23340 13005 24900 13095
rect 23340 12990 23460 13005
rect 24780 12990 24900 13005
rect 25740 13110 25830 13320
rect 25140 13020 25260 13050
rect 25470 12990 25500 13110
rect 25620 12990 25860 13110
rect 26700 12990 26820 13110
rect 22710 12810 22860 12870
rect 22710 12780 22980 12810
rect 22770 12690 22980 12780
rect 25260 12690 25380 12810
rect 18330 12480 18420 12690
rect 19860 12480 19950 12690
rect 20190 12570 20580 12660
rect 20490 12480 20580 12570
rect 22140 12570 22530 12660
rect 22140 12480 22230 12570
rect 22770 12480 22860 12690
rect 25470 12480 25560 12990
rect 25740 12495 25860 12510
rect 26940 12495 27060 13320
rect 29130 13260 29670 13320
rect 28260 13005 29100 13095
rect 29820 13110 29910 13320
rect 30330 13110 30420 13320
rect 30570 13260 31110 13320
rect 29220 13020 29340 13050
rect 29550 12990 29940 13110
rect 30300 12990 30690 13110
rect 31020 13095 31140 13110
rect 31980 13095 32100 13110
rect 31020 13050 32100 13095
rect 30900 13020 32100 13050
rect 31020 13005 32100 13020
rect 31020 12990 31140 13005
rect 31980 12990 32100 13005
rect 25740 12480 27060 12495
rect 16620 12390 16830 12480
rect 16920 12466 17070 12480
rect 16920 12390 16950 12466
rect 16740 12210 16830 12390
rect 16140 11280 16260 11294
rect 16380 11866 16500 11880
rect 16380 11190 16500 11294
rect 16710 11866 16830 11880
rect 16710 11190 16830 11294
rect 16950 11280 17070 11294
rect 17340 12466 17460 12480
rect 17340 11190 17460 11294
rect 17580 12466 17850 12480
rect 17700 12390 17850 12466
rect 18240 12466 18480 12480
rect 17580 11280 17700 11294
rect 17820 12210 17970 12270
rect 17820 11340 17834 12210
rect 17956 11340 17970 12210
rect 17820 11280 17970 11340
rect 18240 11294 18300 12466
rect 18420 11294 18480 12466
rect 18900 12466 19140 12480
rect 18900 12390 19020 12466
rect 18240 11280 18480 11294
rect 18750 12210 18900 12270
rect 18750 11340 18764 12210
rect 18886 11340 18900 12210
rect 17850 11190 17970 11280
rect 18750 11190 18900 11340
rect 19020 11280 19140 11294
rect 19260 12466 19500 12480
rect 19380 12390 19500 12466
rect 19860 12466 20160 12480
rect 19860 12390 19980 12466
rect 19260 11280 19380 11294
rect 19500 12210 19650 12270
rect 19500 11340 19514 12210
rect 19636 11340 19650 12210
rect 19500 11190 19650 11340
rect 19920 11294 19980 12390
rect 20100 11294 20160 12466
rect 20610 12466 20820 12480
rect 20610 12390 20700 12466
rect 19920 11280 20160 11294
rect 20430 12210 20580 12270
rect 20430 11340 20444 12210
rect 20566 11340 20580 12210
rect 20430 11280 20580 11340
rect 20700 11280 20820 11294
rect 21900 12466 22110 12480
rect 22020 12390 22110 12466
rect 22560 12466 22860 12480
rect 21900 11280 22020 11294
rect 22140 12210 22290 12270
rect 22140 11340 22154 12210
rect 22276 11340 22290 12210
rect 22140 11280 22290 11340
rect 22560 11294 22620 12466
rect 22740 12390 22860 12466
rect 22740 11294 22800 12390
rect 23220 12466 23460 12480
rect 23220 12390 23340 12466
rect 22560 11280 22800 11294
rect 23070 12210 23220 12270
rect 23070 11340 23084 12210
rect 23206 11340 23220 12210
rect 20430 11190 20550 11280
rect 22170 11190 22290 11280
rect 23070 11190 23220 11340
rect 23340 11280 23460 11294
rect 25020 12466 25140 12480
rect 25020 11190 25140 11294
rect 25410 12466 25560 12480
rect 25530 12390 25560 12466
rect 25650 12405 27060 12480
rect 25650 12390 25860 12405
rect 25650 12210 25740 12390
rect 25410 11280 25530 11294
rect 25650 11866 25770 11880
rect 25650 11190 25770 11294
rect 26700 11866 26820 11880
rect 26700 11190 26820 11294
rect 26940 11866 27060 12405
rect 27180 12495 27300 12510
rect 27180 12405 27900 12495
rect 27180 12390 27300 12405
rect 29550 12480 29640 12990
rect 29820 12495 29940 12510
rect 29820 12480 30060 12495
rect 29100 12466 29220 12480
rect 26940 11280 27060 11294
rect 27180 11866 27300 11880
rect 27180 11190 27300 11294
rect 29100 11190 29220 11294
rect 29490 12466 29640 12480
rect 29610 12390 29640 12466
rect 29730 12405 30060 12480
rect 29730 12390 29940 12405
rect 30300 12480 30420 12510
rect 30600 12480 30690 12990
rect 30780 12795 30900 12810
rect 30780 12705 31365 12795
rect 30780 12690 30900 12705
rect 31275 12495 31365 12705
rect 31980 12495 32100 12510
rect 30300 12390 30510 12480
rect 30600 12466 30750 12480
rect 30600 12390 30630 12466
rect 29730 12210 29820 12390
rect 30420 12210 30510 12390
rect 29490 11280 29610 11294
rect 29730 11866 29850 11880
rect 29730 11190 29850 11294
rect 30390 11866 30510 11880
rect 30390 11190 30510 11294
rect 30630 11280 30750 11294
rect 31020 12466 31140 12480
rect 31275 12405 32100 12495
rect 31980 12390 32100 12405
rect 31020 11190 31140 11294
rect 31980 11866 32100 11880
rect 31980 11190 32100 11294
rect 32220 11866 32340 13320
rect 32940 13230 33210 13320
rect 32460 12990 32580 13110
rect 32940 12990 33060 13110
rect 33750 13080 33840 13380
rect 34380 13320 34500 13334
rect 34620 13906 34740 13920
rect 34860 13890 34980 14010
rect 34860 13440 34980 13470
rect 35100 13906 35220 13920
rect 34740 13334 35100 13350
rect 34620 13320 35220 13334
rect 35340 13906 35460 13920
rect 35340 13320 35460 13334
rect 36060 13906 36180 14010
rect 36450 13906 36570 13920
rect 36060 13320 36180 13334
rect 36300 13334 36450 13410
rect 36300 13320 36570 13334
rect 37500 13906 37620 14010
rect 37890 13906 38010 13920
rect 37500 13320 37620 13334
rect 37740 13334 37890 13410
rect 37740 13320 38010 13334
rect 38940 13906 39060 14010
rect 39330 13906 39450 13920
rect 38940 13320 39060 13334
rect 39180 13334 39330 13410
rect 39180 13320 39450 13334
rect 40140 13906 40260 13920
rect 40140 13320 40260 13334
rect 40380 13906 40500 13920
rect 40620 13890 40740 14010
rect 40620 13440 40740 13470
rect 40860 13906 40980 13920
rect 40500 13334 40860 13350
rect 40380 13320 40980 13334
rect 41580 13906 41700 13920
rect 41580 13320 41700 13334
rect 41970 13906 42090 14010
rect 42210 13906 42330 13920
rect 42210 13620 42330 13634
rect 43260 13906 43380 14010
rect 42210 13530 42420 13620
rect 41970 13320 42090 13334
rect 34260 13230 34500 13320
rect 34650 13260 35190 13320
rect 33180 13050 33270 13080
rect 33180 12960 33480 13050
rect 33690 12990 33840 13080
rect 33960 13110 34050 13170
rect 34380 12990 34500 13110
rect 34620 13050 34740 13110
rect 35340 13110 35430 13320
rect 34620 13020 34860 13050
rect 34620 12990 34740 13020
rect 35070 12990 35460 13110
rect 36060 13095 36180 13110
rect 35700 13005 36180 13095
rect 36060 12990 36180 13005
rect 33690 12810 33780 12990
rect 33660 12690 33780 12810
rect 34395 12795 34485 12990
rect 34860 12795 34980 12810
rect 34395 12705 34980 12795
rect 34860 12690 34980 12705
rect 33690 12480 33780 12690
rect 35070 12480 35160 12990
rect 35340 12495 35460 12510
rect 36300 12495 36420 13320
rect 36660 13005 37020 13095
rect 37500 13095 37620 13110
rect 37140 13005 37620 13095
rect 37500 12990 37620 13005
rect 35340 12480 36420 12495
rect 32940 12466 33210 12480
rect 32220 11280 32340 11294
rect 32460 11866 32580 11880
rect 32460 11190 32580 11294
rect 33060 12390 33210 12466
rect 33600 12466 33840 12480
rect 32940 11280 33060 11294
rect 33180 12210 33330 12270
rect 33180 11340 33194 12210
rect 33316 11340 33330 12210
rect 33180 11280 33330 11340
rect 33600 11294 33660 12466
rect 33780 11294 33840 12466
rect 34260 12466 34500 12480
rect 34260 12390 34380 12466
rect 33600 11280 33840 11294
rect 34110 12210 34260 12270
rect 34110 11340 34124 12210
rect 34246 11340 34260 12210
rect 33210 11190 33330 11280
rect 34110 11190 34260 11340
rect 34380 11280 34500 11294
rect 34620 12466 34740 12480
rect 34620 11190 34740 11294
rect 35010 12466 35160 12480
rect 35130 12390 35160 12466
rect 35250 12405 36420 12480
rect 35250 12390 35460 12405
rect 35250 12210 35340 12390
rect 35010 11280 35130 11294
rect 35250 11866 35370 11880
rect 35250 11190 35370 11294
rect 36060 11866 36180 11880
rect 36060 11190 36180 11294
rect 36300 11866 36420 12405
rect 36540 12495 36660 12510
rect 37740 12495 37860 13320
rect 38100 13005 38460 13095
rect 38940 13095 39060 13110
rect 38820 13005 39060 13095
rect 38940 12990 39060 13005
rect 39180 12795 39300 13320
rect 40170 13110 40260 13320
rect 40410 13260 40950 13320
rect 41610 13230 41880 13320
rect 41790 13200 41880 13230
rect 40140 13095 40530 13110
rect 40020 13005 40530 13095
rect 41790 13110 42120 13200
rect 40860 13050 40980 13110
rect 40740 13020 40980 13050
rect 40140 12990 40530 13005
rect 40860 12990 40980 13020
rect 41220 13005 41580 13095
rect 39180 12705 39765 12795
rect 36540 12405 37860 12495
rect 36540 12390 36660 12405
rect 36300 11280 36420 11294
rect 36540 11866 36660 11880
rect 36540 11190 36660 11294
rect 37500 11866 37620 11880
rect 37500 11190 37620 11294
rect 37740 11866 37860 12405
rect 37740 11280 37860 11294
rect 37980 11866 38100 11880
rect 37980 11190 38100 11294
rect 38940 11866 39060 11880
rect 38940 11190 39060 11294
rect 39180 11866 39300 12705
rect 39675 12495 39765 12705
rect 40140 12495 40260 12510
rect 39675 12480 40260 12495
rect 40440 12480 40530 12990
rect 40620 12690 40740 12810
rect 41100 12495 41220 12510
rect 41820 12495 42030 12510
rect 39675 12405 40350 12480
rect 40140 12390 40350 12405
rect 40440 12466 40590 12480
rect 40440 12390 40470 12466
rect 40260 12210 40350 12390
rect 39180 11280 39300 11294
rect 39420 11866 39540 11880
rect 39420 11190 39540 11294
rect 40230 11866 40350 11880
rect 40230 11190 40350 11294
rect 40470 11280 40590 11294
rect 40860 12466 40980 12480
rect 41100 12405 42030 12495
rect 41100 12390 41220 12405
rect 41820 12390 42030 12405
rect 42120 12060 42210 13110
rect 42330 12210 42420 13530
rect 43650 13906 43770 13920
rect 43260 13320 43380 13334
rect 43500 13334 43650 13410
rect 43500 13320 43770 13334
rect 44460 13906 44580 13920
rect 44700 13890 44820 14010
rect 44700 13440 44820 13470
rect 44940 13906 45060 13920
rect 44580 13334 44940 13350
rect 44460 13320 45060 13334
rect 45180 13906 45300 13920
rect 45180 13320 45300 13334
rect 46140 13906 46260 14010
rect 46530 13906 46650 13920
rect 46140 13320 46260 13334
rect 46380 13334 46530 13410
rect 46380 13320 46650 13334
rect 47580 13906 47700 13920
rect 47820 13890 47940 14010
rect 47820 13440 47940 13470
rect 48060 13906 48180 13920
rect 47700 13334 48060 13350
rect 47580 13320 48180 13334
rect 48300 13906 48420 13920
rect 48300 13320 48420 13334
rect 49350 13906 49470 13920
rect 49740 13906 49860 14010
rect 49470 13334 49620 13410
rect 49350 13320 49620 13334
rect 49740 13320 49860 13334
rect 43500 12795 43620 13320
rect 44490 13260 45030 13320
rect 44460 13095 44580 13110
rect 44100 13050 44580 13095
rect 45180 13110 45270 13320
rect 44100 13020 44700 13050
rect 44100 13005 44580 13020
rect 44460 12990 44580 13005
rect 44910 12990 45180 13110
rect 45420 13095 45540 13110
rect 46140 13095 46260 13110
rect 45420 13005 46260 13095
rect 45420 12990 45540 13005
rect 46140 12990 46260 13005
rect 44460 12795 44580 12810
rect 43500 12705 44580 12795
rect 42300 12195 42420 12210
rect 42300 12105 43020 12195
rect 42300 12090 42420 12105
rect 41850 11970 42210 12060
rect 41850 11880 41940 11970
rect 42330 11880 42420 12090
rect 40860 11190 40980 11294
rect 41580 11866 41700 11880
rect 41580 11190 41700 11294
rect 41820 11866 41940 11880
rect 41820 11280 41940 11294
rect 42060 11866 42180 11880
rect 42060 11190 42180 11294
rect 42300 11866 42420 11880
rect 42300 11280 42420 11294
rect 43260 11866 43380 11880
rect 43260 11190 43380 11294
rect 43500 11866 43620 12705
rect 44460 12690 44580 12705
rect 44910 12480 45000 12990
rect 45180 12495 45300 12510
rect 46380 12495 46500 13320
rect 47610 13260 48150 13320
rect 46740 13005 47580 13095
rect 48300 13110 48390 13320
rect 47700 13020 47820 13050
rect 48030 12990 48420 13110
rect 46620 12795 46740 12810
rect 46620 12705 47820 12795
rect 46620 12690 46740 12705
rect 45180 12480 46500 12495
rect 44460 12466 44580 12480
rect 43500 11280 43620 11294
rect 43740 11866 43860 11880
rect 43740 11190 43860 11294
rect 44460 11190 44580 11294
rect 44850 12466 45000 12480
rect 44970 12390 45000 12466
rect 45090 12405 46500 12480
rect 45090 12390 45300 12405
rect 45090 12210 45180 12390
rect 44850 11280 44970 11294
rect 45090 11866 45210 11880
rect 45090 11190 45210 11294
rect 46140 11866 46260 11880
rect 46140 11190 46260 11294
rect 46380 11866 46500 12405
rect 46620 12390 46740 12510
rect 48030 12480 48120 12990
rect 49500 12795 49620 13320
rect 49500 12705 49980 12795
rect 48300 12495 48420 12510
rect 48300 12480 49020 12495
rect 47580 12466 47700 12480
rect 46380 11280 46500 11294
rect 46620 11866 46740 11880
rect 46620 11190 46740 11294
rect 47580 11190 47700 11294
rect 47970 12466 48120 12480
rect 48090 12390 48120 12466
rect 48210 12405 49020 12480
rect 48210 12390 48420 12405
rect 49260 12390 49380 12510
rect 48210 12210 48300 12390
rect 47970 11280 48090 11294
rect 48210 11866 48330 11880
rect 48210 11190 48330 11294
rect 49260 11866 49380 11880
rect 49260 11190 49380 11294
rect 49500 11866 49620 12705
rect 49500 11280 49620 11294
rect 49740 11866 49860 11880
rect 49740 11190 49860 11294
rect 1155 11160 54240 11190
rect 1155 11040 1214 11160
rect 2086 11040 5220 11160
rect 5340 11040 5460 11160
rect 5580 11040 5700 11160
rect 5820 11040 5940 11160
rect 6060 11040 6180 11160
rect 6300 11040 6420 11160
rect 6540 11040 6660 11160
rect 6780 11040 6900 11160
rect 7020 11040 7140 11160
rect 7260 11040 7380 11160
rect 7500 11040 7620 11160
rect 7740 11040 7860 11160
rect 7980 11040 8100 11160
rect 8220 11040 8340 11160
rect 8460 11040 8580 11160
rect 8700 11040 8820 11160
rect 8940 11040 9060 11160
rect 9180 11040 9300 11160
rect 9420 11040 9540 11160
rect 9660 11040 9780 11160
rect 9900 11040 10020 11160
rect 10140 11040 10260 11160
rect 10380 11040 10500 11160
rect 10620 11040 10740 11160
rect 10860 11040 10980 11160
rect 11100 11040 11220 11160
rect 11340 11040 11460 11160
rect 11580 11040 11700 11160
rect 11820 11040 11940 11160
rect 12060 11040 12180 11160
rect 12300 11040 12420 11160
rect 12540 11040 12660 11160
rect 12780 11040 12900 11160
rect 13020 11040 13140 11160
rect 13260 11040 13380 11160
rect 13500 11040 13620 11160
rect 13740 11040 13860 11160
rect 13980 11040 14100 11160
rect 14220 11040 14340 11160
rect 14460 11040 14580 11160
rect 14700 11040 14820 11160
rect 14940 11040 15060 11160
rect 15180 11040 15300 11160
rect 15420 11040 15540 11160
rect 15660 11040 15780 11160
rect 15900 11040 16020 11160
rect 16140 11040 16260 11160
rect 16380 11040 16740 11160
rect 16860 11040 16980 11160
rect 17100 11040 17220 11160
rect 17340 11040 17460 11160
rect 17580 11040 17700 11160
rect 17820 11040 17940 11160
rect 18060 11040 18180 11160
rect 18300 11040 18420 11160
rect 18540 11040 18660 11160
rect 18780 11040 18900 11160
rect 19020 11040 19140 11160
rect 19260 11040 19380 11160
rect 19500 11040 19860 11160
rect 19980 11040 20340 11160
rect 20460 11040 20820 11160
rect 20940 11040 21060 11160
rect 21180 11040 21300 11160
rect 21420 11040 21540 11160
rect 21660 11040 21780 11160
rect 21900 11040 22020 11160
rect 22140 11040 22260 11160
rect 22380 11040 22500 11160
rect 22620 11040 22740 11160
rect 22860 11040 22980 11160
rect 23100 11040 23220 11160
rect 23340 11040 23460 11160
rect 23580 11040 23700 11160
rect 23820 11040 23940 11160
rect 24060 11040 24180 11160
rect 24300 11040 24420 11160
rect 24540 11040 24660 11160
rect 24780 11040 24900 11160
rect 25020 11040 25140 11160
rect 25260 11040 25380 11160
rect 25500 11040 25860 11160
rect 25980 11040 26100 11160
rect 26220 11040 26340 11160
rect 26460 11040 26580 11160
rect 26700 11040 26820 11160
rect 26940 11040 27060 11160
rect 27180 11040 27300 11160
rect 27420 11040 27540 11160
rect 27660 11040 27780 11160
rect 27900 11040 28020 11160
rect 28140 11040 28260 11160
rect 28380 11040 28500 11160
rect 28620 11040 28740 11160
rect 28860 11040 28980 11160
rect 29100 11040 29220 11160
rect 29340 11040 29460 11160
rect 29580 11040 29700 11160
rect 29820 11040 29940 11160
rect 30060 11040 30180 11160
rect 30300 11040 30420 11160
rect 30540 11040 30660 11160
rect 30780 11040 30900 11160
rect 31020 11040 31140 11160
rect 31260 11040 31380 11160
rect 31500 11040 31620 11160
rect 31740 11040 31860 11160
rect 31980 11040 32100 11160
rect 32220 11040 32580 11160
rect 32700 11040 32820 11160
rect 32940 11040 33060 11160
rect 33180 11040 33300 11160
rect 33420 11040 33780 11160
rect 33900 11040 34260 11160
rect 34380 11040 34500 11160
rect 34620 11040 34740 11160
rect 34860 11040 34980 11160
rect 35100 11040 35220 11160
rect 35340 11040 35460 11160
rect 35580 11040 35700 11160
rect 35820 11040 35940 11160
rect 36060 11040 36420 11160
rect 36540 11040 36660 11160
rect 36780 11040 36900 11160
rect 37020 11040 37140 11160
rect 37260 11040 37380 11160
rect 37500 11040 37620 11160
rect 37740 11040 37860 11160
rect 37980 11040 38100 11160
rect 38220 11040 38340 11160
rect 38460 11040 38580 11160
rect 38700 11040 38820 11160
rect 38940 11040 39300 11160
rect 39420 11040 39540 11160
rect 39660 11040 39780 11160
rect 39900 11040 40020 11160
rect 40140 11040 40260 11160
rect 40380 11040 40500 11160
rect 40620 11040 40740 11160
rect 40860 11040 40980 11160
rect 41100 11040 41220 11160
rect 41340 11040 41460 11160
rect 41580 11040 41940 11160
rect 42060 11040 42180 11160
rect 42300 11040 42420 11160
rect 42540 11040 42660 11160
rect 42780 11040 42900 11160
rect 43020 11040 43140 11160
rect 43260 11040 43380 11160
rect 43500 11040 43620 11160
rect 43740 11040 43860 11160
rect 43980 11040 44100 11160
rect 44220 11040 44340 11160
rect 44460 11040 44580 11160
rect 44700 11040 44820 11160
rect 44940 11040 45060 11160
rect 45180 11040 45300 11160
rect 45420 11040 45540 11160
rect 45660 11040 45780 11160
rect 45900 11040 46020 11160
rect 46140 11040 46500 11160
rect 46620 11040 46740 11160
rect 46860 11040 46980 11160
rect 47100 11040 47220 11160
rect 47340 11040 47460 11160
rect 47580 11040 47700 11160
rect 47820 11040 47940 11160
rect 48060 11040 48180 11160
rect 48300 11040 48420 11160
rect 48540 11040 48660 11160
rect 48780 11040 48900 11160
rect 49020 11040 49140 11160
rect 49260 11040 49380 11160
rect 49500 11040 49620 11160
rect 49740 11040 49860 11160
rect 49980 11040 50100 11160
rect 50220 11040 53310 11160
rect 54180 11040 54240 11160
rect 1155 11010 54240 11040
rect 5670 10906 5790 11010
rect 5670 10320 5790 10334
rect 5910 10906 6030 10920
rect 5700 9810 5790 9990
rect 5580 9720 5790 9810
rect 5880 9734 5910 9810
rect 5880 9720 6030 9734
rect 6300 10906 6420 11010
rect 6780 10906 6900 11010
rect 6780 10320 6900 10334
rect 7020 10906 7140 10920
rect 6300 9720 6420 9734
rect 6540 9795 6660 9810
rect 7020 9795 7140 10334
rect 7260 10906 7380 11010
rect 8010 10920 8130 11010
rect 7260 10320 7380 10334
rect 7740 10906 7860 10920
rect 5580 9690 5700 9720
rect 5880 9210 5970 9720
rect 6540 9705 7140 9795
rect 6540 9690 6660 9705
rect 6060 9495 6180 9510
rect 6060 9405 6300 9495
rect 6060 9390 6180 9405
rect 5580 9195 5970 9210
rect 5460 9105 5970 9195
rect 6300 9195 6420 9210
rect 6300 9180 6780 9195
rect 5580 9090 5970 9105
rect 6180 9150 6780 9180
rect 5610 8880 5700 9090
rect 6300 9105 6780 9150
rect 6300 9090 6420 9105
rect 5850 8880 6390 8940
rect 7020 8880 7140 9705
rect 7980 10860 8130 10920
rect 7980 9990 7994 10860
rect 8116 9990 8130 10860
rect 7980 9930 8130 9990
rect 8400 10906 8640 10920
rect 7860 9734 8010 9810
rect 7740 9720 8010 9734
rect 8400 9734 8460 10906
rect 8580 9734 8640 10906
rect 8910 10860 9060 11010
rect 8910 9990 8924 10860
rect 9046 9990 9060 10860
rect 8910 9930 9060 9990
rect 9180 10906 9300 10920
rect 8400 9720 8640 9734
rect 9060 9734 9180 9810
rect 9660 10906 9780 10920
rect 9540 10605 9660 10695
rect 9060 9720 9300 9734
rect 9660 10320 9780 10334
rect 9900 10906 10020 11010
rect 9900 10320 10020 10334
rect 10140 10906 10260 10920
rect 10140 10320 10260 10334
rect 10380 10906 10500 11010
rect 10380 10320 10500 10334
rect 11340 10906 11460 11010
rect 11340 10320 11460 10334
rect 11580 10906 11700 10920
rect 9660 10110 9750 10320
rect 10140 10230 10230 10320
rect 9870 10140 10230 10230
rect 9660 9990 9780 10110
rect 8490 9510 8580 9720
rect 8460 9390 8580 9510
rect 7740 9090 7860 9210
rect 7980 9150 8280 9240
rect 8490 9210 8580 9390
rect 7980 9120 8070 9150
rect 8490 9120 8640 9210
rect 7740 8880 8010 8970
rect 5580 8866 5700 8880
rect 5580 8280 5700 8294
rect 5820 8866 6420 8880
rect 5940 8850 6300 8866
rect 5820 8280 5940 8294
rect 6060 8730 6180 8760
rect 6060 8190 6180 8310
rect 6300 8280 6420 8294
rect 6780 8866 6900 8880
rect 7020 8866 7290 8880
rect 7020 8790 7170 8866
rect 6780 8190 6900 8294
rect 7170 8280 7290 8294
rect 7740 8866 7860 8880
rect 8550 8820 8640 9120
rect 9180 9195 9300 9210
rect 9180 9105 9420 9195
rect 9180 9090 9300 9105
rect 8760 9030 8850 9090
rect 9060 8880 9300 8970
rect 7740 8280 7860 8294
rect 7980 8746 8130 8790
rect 7980 8324 7994 8746
rect 8116 8324 8130 8746
rect 7980 8280 8130 8324
rect 8400 8760 8640 8820
rect 9180 8866 9300 8880
rect 8400 8340 8460 8760
rect 8580 8340 8640 8760
rect 8400 8280 8640 8340
rect 8910 8746 9060 8790
rect 8910 8324 8924 8746
rect 9046 8324 9060 8746
rect 8010 8190 8130 8280
rect 8910 8190 9060 8324
rect 9660 8670 9750 9990
rect 9870 9090 9960 10140
rect 10050 9690 10140 9810
rect 11340 9795 11460 9810
rect 11220 9705 11460 9795
rect 11340 9690 11460 9705
rect 9960 9000 10290 9090
rect 10200 8970 10290 9000
rect 10200 8880 10470 8970
rect 11580 8880 11700 10334
rect 11820 10906 11940 11010
rect 14010 10920 14130 11010
rect 11820 10320 11940 10334
rect 13740 10906 13860 10920
rect 13980 10860 14130 10920
rect 13980 9990 13994 10860
rect 14116 9990 14130 10860
rect 13980 9930 14130 9990
rect 14400 10906 14640 10920
rect 13860 9734 14010 9810
rect 13740 9720 14010 9734
rect 14400 9734 14460 10906
rect 14580 9734 14640 10906
rect 14910 10860 15060 11010
rect 14910 9990 14924 10860
rect 15046 9990 15060 10860
rect 14910 9930 15060 9990
rect 15180 10906 15300 10920
rect 14400 9720 14640 9734
rect 15060 9734 15180 9810
rect 16380 10906 16500 11010
rect 16380 10320 16500 10334
rect 16620 10906 16740 10920
rect 15060 9720 15300 9734
rect 14490 9510 14580 9720
rect 14460 9495 14580 9510
rect 16380 9495 16500 9510
rect 14460 9405 16500 9495
rect 14460 9390 14580 9405
rect 16380 9390 16500 9405
rect 11820 9195 11940 9210
rect 11820 9105 12540 9195
rect 11820 9090 11940 9105
rect 13740 9195 13860 9210
rect 12900 9105 13860 9195
rect 13740 9090 13860 9105
rect 13980 9150 14280 9240
rect 14490 9210 14580 9390
rect 13980 9120 14070 9150
rect 14490 9120 14640 9210
rect 13740 8880 14010 8970
rect 9990 8866 10110 8880
rect 9660 8580 9870 8670
rect 9180 8280 9300 8294
rect 9750 8566 9870 8580
rect 9750 8280 9870 8294
rect 9990 8190 10110 8294
rect 10380 8866 10500 8880
rect 10380 8280 10500 8294
rect 11430 8866 11700 8880
rect 11550 8790 11700 8866
rect 11820 8866 11940 8880
rect 11430 8280 11550 8294
rect 11820 8190 11940 8294
rect 13740 8866 13860 8880
rect 14550 8820 14640 9120
rect 16380 9090 16500 9210
rect 14760 9030 14850 9090
rect 15060 8880 15300 8970
rect 16620 8880 16740 10334
rect 16860 10906 16980 11010
rect 17610 10920 17730 11010
rect 16860 10320 16980 10334
rect 17340 10906 17460 10920
rect 16860 9795 16980 9810
rect 16860 9705 17100 9795
rect 16860 9690 16980 9705
rect 17580 10860 17730 10920
rect 17580 9990 17594 10860
rect 17716 9990 17730 10860
rect 17580 9930 17730 9990
rect 18000 10906 18240 10920
rect 17460 9734 17550 9810
rect 17340 9720 17550 9734
rect 18000 9734 18060 10906
rect 18180 9810 18240 10906
rect 18510 10860 18660 11010
rect 18510 9990 18524 10860
rect 18646 9990 18660 10860
rect 18510 9930 18660 9990
rect 18780 10906 18900 10920
rect 18180 9734 18300 9810
rect 18000 9720 18300 9734
rect 18660 9734 18780 9810
rect 18660 9720 18900 9734
rect 19260 10906 19380 10920
rect 19500 10860 19650 11010
rect 20430 10920 20550 11010
rect 19500 9990 19514 10860
rect 19636 9990 19650 10860
rect 19500 9930 19650 9990
rect 19920 10906 20160 10920
rect 19380 9734 19500 9810
rect 19260 9720 19500 9734
rect 19920 9734 19980 10906
rect 20100 9734 20160 10906
rect 20430 10860 20580 10920
rect 20430 9990 20444 10860
rect 20566 9990 20580 10860
rect 20430 9930 20580 9990
rect 20700 10906 20820 10920
rect 19920 9720 20160 9734
rect 20550 9734 20700 9810
rect 21180 10906 21300 11010
rect 21180 10320 21300 10334
rect 21420 10906 21540 10920
rect 20550 9720 20820 9734
rect 17580 9630 17670 9720
rect 17580 9540 17970 9630
rect 18210 9510 18300 9720
rect 19980 9510 20070 9720
rect 21180 9795 21300 9810
rect 21060 9705 21300 9795
rect 21180 9690 21300 9705
rect 18210 9420 18420 9510
rect 19980 9495 20100 9510
rect 17760 9330 18030 9420
rect 17940 9240 18030 9330
rect 18150 9390 18420 9420
rect 19035 9405 20100 9495
rect 18150 9330 18300 9390
rect 17340 9090 17460 9210
rect 17580 9090 17850 9180
rect 17760 9030 17850 9090
rect 17340 8880 17550 8970
rect 17760 8940 17820 9030
rect 13740 8280 13860 8294
rect 13980 8746 14130 8790
rect 13980 8324 13994 8746
rect 14116 8324 14130 8746
rect 13980 8280 14130 8324
rect 14400 8760 14640 8820
rect 15180 8866 15300 8880
rect 14400 8340 14460 8760
rect 14580 8340 14640 8760
rect 14400 8280 14640 8340
rect 14910 8746 15060 8790
rect 14910 8324 14924 8746
rect 15046 8324 15060 8746
rect 14010 8190 14130 8280
rect 14910 8190 15060 8324
rect 15180 8280 15300 8294
rect 16380 8866 16500 8880
rect 16620 8866 16890 8880
rect 16620 8790 16770 8866
rect 16380 8190 16500 8294
rect 16770 8280 16890 8294
rect 17340 8866 17460 8880
rect 18150 8820 18240 9330
rect 18780 9195 18900 9210
rect 19035 9195 19125 9405
rect 19980 9390 20100 9405
rect 19980 9210 20070 9390
rect 18780 9105 19125 9195
rect 18780 9090 18900 9105
rect 19260 9090 19380 9210
rect 18360 9030 18450 9090
rect 19710 9030 19800 9090
rect 19920 9120 20070 9210
rect 20280 9150 20580 9240
rect 20490 9120 20580 9150
rect 18660 8880 18900 8970
rect 17340 8280 17460 8294
rect 17580 8746 17730 8790
rect 17580 8324 17594 8746
rect 17716 8324 17730 8746
rect 17580 8280 17730 8324
rect 18000 8760 18240 8820
rect 18780 8866 18900 8880
rect 18000 8340 18060 8760
rect 18180 8340 18240 8760
rect 18000 8280 18240 8340
rect 18510 8746 18660 8790
rect 18510 8324 18524 8746
rect 18646 8324 18660 8746
rect 17610 8190 17730 8280
rect 18510 8190 18660 8324
rect 18780 8280 18900 8294
rect 19260 8880 19500 8970
rect 19260 8866 19380 8880
rect 19920 8820 20010 9120
rect 20820 9105 21180 9195
rect 20550 8880 20820 8970
rect 21420 8910 21540 10334
rect 21660 10906 21780 11010
rect 21660 10320 21780 10334
rect 21900 10906 22020 10920
rect 22140 10860 22290 11010
rect 23070 10920 23190 11010
rect 22140 9990 22154 10860
rect 22276 9990 22290 10860
rect 22140 9930 22290 9990
rect 22560 10906 22800 10920
rect 22020 9734 22140 9810
rect 21900 9720 22140 9734
rect 22560 9734 22620 10906
rect 22740 9734 22800 10906
rect 23070 10860 23220 10920
rect 23070 9990 23084 10860
rect 23206 9990 23220 10860
rect 23070 9930 23220 9990
rect 23340 10906 23460 10920
rect 22560 9720 22800 9734
rect 23190 9734 23340 9810
rect 23820 10906 23940 11010
rect 23820 10320 23940 10334
rect 24060 10906 24180 10920
rect 23190 9720 23460 9734
rect 22620 9510 22710 9720
rect 22620 9390 22740 9510
rect 22620 9210 22710 9390
rect 21660 9090 21780 9210
rect 22350 9030 22440 9090
rect 22560 9120 22710 9210
rect 22920 9150 23220 9240
rect 23130 9120 23220 9150
rect 20700 8866 20820 8880
rect 19260 8280 19380 8294
rect 19500 8746 19650 8790
rect 19500 8324 19514 8746
rect 19636 8324 19650 8746
rect 19500 8190 19650 8324
rect 19920 8760 20160 8820
rect 19920 8340 19980 8760
rect 20100 8340 20160 8760
rect 19920 8280 20160 8340
rect 20430 8746 20580 8790
rect 20430 8324 20444 8746
rect 20566 8324 20580 8746
rect 20430 8280 20580 8324
rect 20700 8280 20820 8294
rect 21270 8866 21420 8880
rect 21390 8790 21420 8866
rect 21900 8880 22140 8970
rect 21660 8866 21780 8880
rect 21270 8280 21390 8294
rect 20430 8190 20550 8280
rect 21660 8190 21780 8294
rect 21900 8866 22020 8880
rect 22560 8820 22650 9120
rect 23190 8880 23460 8970
rect 24060 8880 24180 10334
rect 24300 10906 24420 11010
rect 25770 10920 25890 11010
rect 24300 10320 24420 10334
rect 25500 10906 25620 10920
rect 24300 9795 24420 9810
rect 24300 9705 24540 9795
rect 24300 9690 24420 9705
rect 24660 9705 25260 9795
rect 25740 10860 25890 10920
rect 25740 9990 25754 10860
rect 25876 9990 25890 10860
rect 25740 9930 25890 9990
rect 26160 10906 26400 10920
rect 25620 9734 25770 9810
rect 25500 9720 25770 9734
rect 26160 9734 26220 10906
rect 26340 9734 26400 10906
rect 26670 10860 26820 11010
rect 26670 9990 26684 10860
rect 26806 9990 26820 10860
rect 26670 9930 26820 9990
rect 26940 10906 27060 10920
rect 26160 9720 26400 9734
rect 26820 9734 26940 9810
rect 27900 10906 28020 11010
rect 27900 10320 28020 10334
rect 28140 10906 28260 10920
rect 26820 9720 27060 9734
rect 26250 9510 26340 9720
rect 26220 9390 26340 9510
rect 24420 9105 25020 9195
rect 25500 9195 25620 9210
rect 25140 9105 25620 9195
rect 25500 9090 25620 9105
rect 25740 9150 26040 9240
rect 26250 9210 26340 9390
rect 25740 9120 25830 9150
rect 26250 9120 26400 9210
rect 25500 8880 25770 8970
rect 23340 8866 23460 8880
rect 21900 8280 22020 8294
rect 22140 8746 22290 8790
rect 22140 8324 22154 8746
rect 22276 8324 22290 8746
rect 22140 8190 22290 8324
rect 22560 8760 22800 8820
rect 22560 8340 22620 8760
rect 22740 8340 22800 8760
rect 22560 8280 22800 8340
rect 23070 8746 23220 8790
rect 23070 8324 23084 8746
rect 23206 8324 23220 8746
rect 23070 8280 23220 8324
rect 23340 8280 23460 8294
rect 23820 8866 23940 8880
rect 24060 8866 24330 8880
rect 24060 8790 24210 8866
rect 23070 8190 23190 8280
rect 23820 8190 23940 8294
rect 24210 8280 24330 8294
rect 25500 8866 25620 8880
rect 26310 8820 26400 9120
rect 27900 9195 28020 9210
rect 27540 9105 28020 9195
rect 27900 9090 28020 9105
rect 26520 9030 26610 9090
rect 26820 8880 27060 8970
rect 28140 8895 28260 10334
rect 28380 10906 28500 11010
rect 28380 10320 28500 10334
rect 29340 10890 29460 10920
rect 29580 10890 29700 11010
rect 30540 10890 30660 11010
rect 30780 10890 30900 10920
rect 28500 9705 28860 9795
rect 29100 8895 29220 8910
rect 25500 8280 25620 8294
rect 25740 8746 25890 8790
rect 25740 8324 25754 8746
rect 25876 8324 25890 8746
rect 25740 8280 25890 8324
rect 26160 8760 26400 8820
rect 26940 8866 27060 8880
rect 26160 8340 26220 8760
rect 26340 8340 26400 8760
rect 26160 8280 26400 8340
rect 26670 8746 26820 8790
rect 26670 8324 26684 8746
rect 26806 8324 26820 8746
rect 25770 8190 25890 8280
rect 26670 8190 26820 8324
rect 26940 8280 27060 8294
rect 27900 8866 28020 8880
rect 28140 8866 29220 8895
rect 28140 8790 28290 8866
rect 27900 8190 28020 8294
rect 28410 8805 29220 8866
rect 29100 8790 29220 8805
rect 28290 8280 28410 8294
rect 29340 8550 29460 10320
rect 30780 9495 30900 10320
rect 31740 10906 31860 11010
rect 31740 9720 31860 9734
rect 32130 10906 32250 10920
rect 32370 10906 32490 11010
rect 32370 10320 32490 10334
rect 33180 10906 33300 10920
rect 32250 9734 32280 9810
rect 32130 9720 32280 9734
rect 32370 9720 32460 9990
rect 31980 9495 32100 9510
rect 30780 9405 32100 9495
rect 29820 8895 29940 8910
rect 30540 8895 30660 8910
rect 29820 8805 30660 8895
rect 29820 8790 29940 8805
rect 30540 8790 30660 8805
rect 29580 8550 29700 8580
rect 29580 8190 29700 8280
rect 30540 8550 30660 8580
rect 30780 8550 30900 9405
rect 31980 9390 32100 9405
rect 32190 9210 32280 9720
rect 33420 10860 33570 11010
rect 34350 10920 34470 11010
rect 33420 9990 33434 10860
rect 33556 9990 33570 10860
rect 33420 9930 33570 9990
rect 33840 10906 34080 10920
rect 33300 9734 33420 9810
rect 33180 9720 33420 9734
rect 33840 9810 33900 10906
rect 33780 9734 33900 9810
rect 34020 9734 34080 10906
rect 34350 10860 34500 10920
rect 34350 9990 34364 10860
rect 34486 9990 34500 10860
rect 34350 9930 34500 9990
rect 34620 10906 34740 10920
rect 33780 9720 34080 9734
rect 34530 9734 34620 9810
rect 34530 9720 34740 9734
rect 35580 10906 35700 10920
rect 35580 10320 35700 10334
rect 35820 10906 35940 11010
rect 35820 10320 35940 10334
rect 36060 10906 36180 10920
rect 36060 10320 36180 10334
rect 36300 10906 36420 11010
rect 36300 10320 36420 10334
rect 36780 10906 36900 11010
rect 36780 10320 36900 10334
rect 37020 10906 37140 10920
rect 35580 10110 35670 10320
rect 36060 10230 36150 10320
rect 35790 10140 36150 10230
rect 33780 9510 33870 9720
rect 34410 9630 34500 9720
rect 34110 9540 34500 9630
rect 33660 9420 33870 9510
rect 33660 9390 33930 9420
rect 33780 9330 33930 9390
rect 31020 9195 31140 9210
rect 31020 9105 31740 9195
rect 31020 9090 31140 9105
rect 31860 9150 31980 9180
rect 32190 9090 32220 9210
rect 32340 9090 32580 9210
rect 31770 8880 32310 8940
rect 32460 8880 32550 9090
rect 33630 9030 33720 9090
rect 33180 8880 33420 8970
rect 31740 8866 32340 8880
rect 31860 8850 32220 8866
rect 31740 8280 31860 8294
rect 31980 8730 32100 8760
rect 30540 8190 30660 8280
rect 31980 8190 32100 8310
rect 32220 8280 32340 8294
rect 32460 8866 32580 8880
rect 32460 8280 32580 8294
rect 33180 8866 33300 8880
rect 33840 8820 33930 9330
rect 34050 9330 34320 9420
rect 34050 9240 34140 9330
rect 34230 9090 34500 9180
rect 34620 9195 34740 9210
rect 34620 9105 35340 9195
rect 34620 9090 34740 9105
rect 34230 9030 34320 9090
rect 34260 8940 34320 9030
rect 34530 8880 34740 8970
rect 34620 8866 34740 8880
rect 33180 8280 33300 8294
rect 33420 8746 33570 8790
rect 33420 8324 33434 8746
rect 33556 8324 33570 8746
rect 33420 8190 33570 8324
rect 33840 8760 34080 8820
rect 33840 8340 33900 8760
rect 34020 8340 34080 8760
rect 33840 8280 34080 8340
rect 34350 8746 34500 8790
rect 34350 8324 34364 8746
rect 34486 8324 34500 8746
rect 34350 8280 34500 8324
rect 35580 8670 35670 9990
rect 35790 9090 35880 10140
rect 35970 9795 36180 9810
rect 36780 9795 36900 9810
rect 35970 9705 36900 9795
rect 35970 9690 36180 9705
rect 36780 9690 36900 9705
rect 36780 9195 36900 9210
rect 36420 9105 36900 9195
rect 36780 9090 36900 9105
rect 35880 9000 36210 9090
rect 36120 8970 36210 9000
rect 36120 8880 36390 8970
rect 37020 8880 37140 10334
rect 37260 10906 37380 11010
rect 37260 10320 37380 10334
rect 37740 10906 37860 10920
rect 37740 10320 37860 10334
rect 37980 10906 38100 11010
rect 37980 10320 38100 10334
rect 38220 10906 38340 10920
rect 38220 10320 38340 10334
rect 38460 10906 38580 11010
rect 38460 10320 38580 10334
rect 38940 10906 39060 11010
rect 37740 10110 37830 10320
rect 38220 10230 38310 10320
rect 37950 10140 38310 10230
rect 37740 9990 37860 10110
rect 35910 8866 36030 8880
rect 35580 8580 35790 8670
rect 34620 8280 34740 8294
rect 35670 8566 35790 8580
rect 35670 8280 35790 8294
rect 34350 8190 34470 8280
rect 35910 8190 36030 8294
rect 36300 8866 36420 8880
rect 36300 8280 36420 8294
rect 36780 8866 36900 8880
rect 37020 8866 37290 8880
rect 37020 8790 37170 8866
rect 36780 8190 36900 8294
rect 37740 8670 37830 9990
rect 37950 9090 38040 10140
rect 38130 9690 38340 9810
rect 38940 9720 39060 9734
rect 39330 10906 39450 10920
rect 39570 10906 39690 11010
rect 39570 10320 39690 10334
rect 40380 10906 40500 11010
rect 40380 10320 40500 10334
rect 40620 10906 40740 10920
rect 39570 9810 39660 9990
rect 39450 9734 39480 9810
rect 39330 9720 39480 9734
rect 39570 9795 39780 9810
rect 40620 9795 40740 10334
rect 40860 10906 40980 11010
rect 40860 10320 40980 10334
rect 41580 10906 41700 11010
rect 41580 10320 41700 10334
rect 41820 10906 41940 10920
rect 39570 9720 40740 9795
rect 39180 9390 39300 9510
rect 39390 9210 39480 9720
rect 39660 9705 40740 9720
rect 39660 9690 39780 9705
rect 39060 9150 39180 9180
rect 38040 9000 38370 9090
rect 39390 9090 39780 9210
rect 40380 9195 40500 9210
rect 40020 9105 40500 9195
rect 40380 9090 40500 9105
rect 38280 8970 38370 9000
rect 38280 8880 38550 8970
rect 38970 8880 39510 8940
rect 39660 8880 39750 9090
rect 40620 8880 40740 9705
rect 41580 9195 41700 9210
rect 41220 9105 41700 9195
rect 41580 9090 41700 9105
rect 41820 9195 41940 10334
rect 42060 10906 42180 11010
rect 42810 10920 42930 11010
rect 42060 10320 42180 10334
rect 42540 10906 42660 10920
rect 42060 9690 42180 9810
rect 42780 10860 42930 10920
rect 42780 9990 42794 10860
rect 42916 9990 42930 10860
rect 42780 9930 42930 9990
rect 43200 10906 43440 10920
rect 42660 9734 42810 9810
rect 42540 9720 42810 9734
rect 43200 9734 43260 10906
rect 43380 9734 43440 10906
rect 43710 10860 43860 11010
rect 45450 10920 45570 11010
rect 43710 9990 43724 10860
rect 43846 9990 43860 10860
rect 43710 9930 43860 9990
rect 43980 10906 44100 10920
rect 43200 9720 43440 9734
rect 43860 9734 43980 9810
rect 43860 9720 44100 9734
rect 45180 10906 45300 10920
rect 45420 10860 45570 10920
rect 45420 9990 45434 10860
rect 45556 9990 45570 10860
rect 45420 9930 45570 9990
rect 45840 10906 46080 10920
rect 45300 9734 45450 9810
rect 45180 9720 45450 9734
rect 45840 9734 45900 10906
rect 46020 9734 46080 10906
rect 46350 10860 46500 11010
rect 46350 9990 46364 10860
rect 46486 9990 46500 10860
rect 46350 9930 46500 9990
rect 46620 10906 46740 10920
rect 45840 9720 46080 9734
rect 46500 9734 46620 9810
rect 47580 10906 47700 11010
rect 47580 10320 47700 10334
rect 47820 10906 47940 10920
rect 46500 9720 46740 9734
rect 43290 9510 43380 9720
rect 43260 9390 43380 9510
rect 44100 9405 44460 9495
rect 45930 9510 46020 9720
rect 47820 9795 47940 10334
rect 48060 10906 48180 11010
rect 48060 10320 48180 10334
rect 49020 10906 49140 11010
rect 49020 10320 49140 10334
rect 49260 10906 49380 10920
rect 49020 9795 49140 9810
rect 47820 9705 49140 9795
rect 45900 9495 46020 9510
rect 45900 9405 47580 9495
rect 45900 9390 46020 9405
rect 42300 9195 42420 9210
rect 41820 9105 42420 9195
rect 41820 8880 41940 9105
rect 42300 9090 42420 9105
rect 42780 9150 43080 9240
rect 43290 9210 43380 9390
rect 42780 9120 42870 9150
rect 43290 9120 43440 9210
rect 42540 8880 42810 8970
rect 38070 8866 38190 8880
rect 37740 8580 37950 8670
rect 37170 8280 37290 8294
rect 37830 8566 37950 8580
rect 37830 8280 37950 8294
rect 38070 8190 38190 8294
rect 38460 8866 38580 8880
rect 38460 8280 38580 8294
rect 38940 8866 39540 8880
rect 39060 8850 39420 8866
rect 38940 8280 39060 8294
rect 39180 8730 39300 8760
rect 39180 8190 39300 8310
rect 39420 8280 39540 8294
rect 39660 8866 39780 8880
rect 39660 8280 39780 8294
rect 40380 8866 40500 8880
rect 40620 8866 40890 8880
rect 40620 8790 40770 8866
rect 40380 8190 40500 8294
rect 40770 8280 40890 8294
rect 41580 8866 41700 8880
rect 41820 8866 42090 8880
rect 41820 8790 41970 8866
rect 41580 8190 41700 8294
rect 41970 8280 42090 8294
rect 42540 8866 42660 8880
rect 43350 8820 43440 9120
rect 43980 9090 44100 9210
rect 45420 9150 45720 9240
rect 45930 9210 46020 9390
rect 45420 9120 45510 9150
rect 45930 9120 46080 9210
rect 43560 9030 43650 9090
rect 43860 8880 44100 8970
rect 42540 8280 42660 8294
rect 42780 8746 42930 8790
rect 42780 8324 42794 8746
rect 42916 8324 42930 8746
rect 42780 8280 42930 8324
rect 43200 8760 43440 8820
rect 43980 8866 44100 8880
rect 43200 8340 43260 8760
rect 43380 8340 43440 8760
rect 43200 8280 43440 8340
rect 43710 8746 43860 8790
rect 43710 8324 43724 8746
rect 43846 8324 43860 8746
rect 42810 8190 42930 8280
rect 43710 8190 43860 8324
rect 43980 8280 44100 8294
rect 45180 8880 45450 8970
rect 45180 8866 45300 8880
rect 45990 8820 46080 9120
rect 46620 9195 46740 9210
rect 46620 9105 46860 9195
rect 46620 9090 46740 9105
rect 46200 9030 46290 9090
rect 46500 8880 46740 8970
rect 47820 8880 47940 9705
rect 49020 9690 49140 9705
rect 48060 9195 48180 9210
rect 48060 9105 48300 9195
rect 48060 9090 48180 9105
rect 49260 8880 49380 10334
rect 49500 10906 49620 11010
rect 49500 10320 49620 10334
rect 49500 9090 49620 9210
rect 45180 8280 45300 8294
rect 45420 8746 45570 8790
rect 45420 8324 45434 8746
rect 45556 8324 45570 8746
rect 45420 8280 45570 8324
rect 45840 8760 46080 8820
rect 46620 8866 46740 8880
rect 45840 8340 45900 8760
rect 46020 8340 46080 8760
rect 45840 8280 46080 8340
rect 46350 8746 46500 8790
rect 46350 8324 46364 8746
rect 46486 8324 46500 8746
rect 45450 8190 45570 8280
rect 46350 8190 46500 8324
rect 46620 8280 46740 8294
rect 47670 8866 47940 8880
rect 47790 8790 47940 8866
rect 48060 8866 48180 8880
rect 47670 8280 47790 8294
rect 48060 8190 48180 8294
rect 49110 8866 49380 8880
rect 49230 8790 49380 8866
rect 49500 8866 49620 8880
rect 49110 8280 49230 8294
rect 49500 8190 49620 8294
rect 3135 8160 52260 8190
rect 3135 8040 3194 8160
rect 4066 8040 5220 8160
rect 5340 8040 5460 8160
rect 5580 8040 5700 8160
rect 5820 8040 5940 8160
rect 6060 8040 6180 8160
rect 6300 8040 6420 8160
rect 6540 8040 6660 8160
rect 6780 8040 7140 8160
rect 7260 8040 7380 8160
rect 7500 8040 7620 8160
rect 7740 8040 7860 8160
rect 7980 8040 8100 8160
rect 8220 8040 8340 8160
rect 8460 8040 8580 8160
rect 8700 8040 9060 8160
rect 9180 8040 9300 8160
rect 9420 8040 9540 8160
rect 9660 8040 9780 8160
rect 9900 8040 10020 8160
rect 10140 8040 10260 8160
rect 10380 8040 10500 8160
rect 10620 8040 10740 8160
rect 10860 8040 10980 8160
rect 11100 8040 11220 8160
rect 11340 8040 11460 8160
rect 11580 8040 11700 8160
rect 11820 8040 11940 8160
rect 12060 8040 12180 8160
rect 12300 8040 12420 8160
rect 12540 8040 12660 8160
rect 12780 8040 12900 8160
rect 13020 8040 13140 8160
rect 13260 8040 13380 8160
rect 13500 8040 13620 8160
rect 13740 8040 14100 8160
rect 14220 8040 14580 8160
rect 14700 8040 14820 8160
rect 14940 8040 15060 8160
rect 15180 8040 15300 8160
rect 15420 8040 15540 8160
rect 15660 8040 15780 8160
rect 15900 8040 16020 8160
rect 16140 8040 16260 8160
rect 16380 8040 16500 8160
rect 16620 8040 16740 8160
rect 16860 8040 16980 8160
rect 17100 8040 17220 8160
rect 17340 8040 17460 8160
rect 17580 8040 17700 8160
rect 17820 8040 17940 8160
rect 18060 8040 18180 8160
rect 18300 8040 18420 8160
rect 18540 8040 18660 8160
rect 18780 8040 18900 8160
rect 19020 8040 19140 8160
rect 19260 8040 19380 8160
rect 19500 8040 19620 8160
rect 19740 8040 19860 8160
rect 19980 8040 20100 8160
rect 20220 8040 20340 8160
rect 20460 8040 20580 8160
rect 20700 8040 20820 8160
rect 20940 8040 21060 8160
rect 21180 8040 21300 8160
rect 21420 8040 21540 8160
rect 21660 8040 21780 8160
rect 21900 8040 22020 8160
rect 22140 8040 22260 8160
rect 22380 8040 22500 8160
rect 22620 8040 22740 8160
rect 22860 8040 22980 8160
rect 23100 8040 23220 8160
rect 23340 8040 23460 8160
rect 23580 8040 23700 8160
rect 23820 8040 23940 8160
rect 24060 8040 24180 8160
rect 24300 8040 24420 8160
rect 24540 8040 24660 8160
rect 24780 8040 24900 8160
rect 25020 8040 25140 8160
rect 25260 8040 25380 8160
rect 25500 8040 25620 8160
rect 25740 8040 25860 8160
rect 25980 8040 26100 8160
rect 26220 8040 26340 8160
rect 26460 8040 26580 8160
rect 26700 8040 26820 8160
rect 26940 8040 27060 8160
rect 27180 8040 27300 8160
rect 27420 8040 27540 8160
rect 27660 8040 27780 8160
rect 27900 8040 28260 8160
rect 28380 8040 28500 8160
rect 28620 8040 28740 8160
rect 28860 8040 28980 8160
rect 29100 8040 29220 8160
rect 29340 8040 29460 8160
rect 29580 8040 29700 8160
rect 29820 8040 29940 8160
rect 30060 8040 30180 8160
rect 30300 8040 30420 8160
rect 30540 8040 30900 8160
rect 31020 8040 31140 8160
rect 31260 8040 31380 8160
rect 31500 8040 31620 8160
rect 31740 8040 31860 8160
rect 31980 8040 32100 8160
rect 32220 8040 32340 8160
rect 32460 8040 32580 8160
rect 32700 8040 32820 8160
rect 32940 8040 33060 8160
rect 33180 8040 33300 8160
rect 33420 8040 33540 8160
rect 33660 8040 33780 8160
rect 33900 8040 34020 8160
rect 34140 8040 34260 8160
rect 34380 8040 34500 8160
rect 34620 8040 34740 8160
rect 34860 8040 34980 8160
rect 35100 8040 35220 8160
rect 35340 8040 35460 8160
rect 35580 8040 35700 8160
rect 35820 8040 35940 8160
rect 36060 8040 36420 8160
rect 36540 8040 36660 8160
rect 36780 8040 36900 8160
rect 37020 8040 37140 8160
rect 37260 8040 37380 8160
rect 37500 8040 37620 8160
rect 37740 8040 37860 8160
rect 37980 8040 38100 8160
rect 38220 8040 38340 8160
rect 38460 8040 38580 8160
rect 38700 8040 38820 8160
rect 38940 8040 39300 8160
rect 39420 8040 39540 8160
rect 39660 8040 39780 8160
rect 39900 8040 40020 8160
rect 40140 8040 40260 8160
rect 40380 8040 40740 8160
rect 40860 8040 40980 8160
rect 41100 8040 41220 8160
rect 41340 8040 41460 8160
rect 41580 8040 41700 8160
rect 41820 8040 41940 8160
rect 42060 8040 42180 8160
rect 42300 8040 42420 8160
rect 42540 8040 42660 8160
rect 42780 8040 42900 8160
rect 43020 8040 43140 8160
rect 43260 8040 43380 8160
rect 43500 8040 43620 8160
rect 43740 8040 43860 8160
rect 43980 8040 44100 8160
rect 44220 8040 44340 8160
rect 44460 8040 44580 8160
rect 44700 8040 44820 8160
rect 44940 8040 45060 8160
rect 45180 8040 45300 8160
rect 45420 8040 45540 8160
rect 45660 8040 45780 8160
rect 45900 8040 46020 8160
rect 46140 8040 46260 8160
rect 46380 8040 46500 8160
rect 46620 8040 46740 8160
rect 46860 8040 46980 8160
rect 47100 8040 47220 8160
rect 47340 8040 47460 8160
rect 47580 8040 47700 8160
rect 47820 8040 48180 8160
rect 48300 8040 48420 8160
rect 48540 8040 48660 8160
rect 48780 8040 48900 8160
rect 49020 8040 49140 8160
rect 49260 8040 49380 8160
rect 49500 8040 49620 8160
rect 49740 8040 49860 8160
rect 49980 8040 50100 8160
rect 50220 8040 51330 8160
rect 52200 8040 52260 8160
rect 3135 8010 52260 8040
rect 5580 7906 5700 7920
rect 5820 7876 5970 8010
rect 6750 7920 6870 8010
rect 8220 7920 8340 8010
rect 5820 7454 5834 7876
rect 5956 7454 5970 7876
rect 5820 7410 5970 7454
rect 6240 7860 6480 7920
rect 6240 7440 6300 7860
rect 6420 7440 6480 7860
rect 5580 7320 5700 7334
rect 6240 7380 6480 7440
rect 6750 7876 6900 7920
rect 6750 7454 6764 7876
rect 6886 7454 6900 7876
rect 6750 7410 6900 7454
rect 7020 7906 7140 7920
rect 5580 7230 5820 7320
rect 6030 7110 6120 7170
rect 5580 6990 5700 7110
rect 6240 7080 6330 7380
rect 7380 7650 7980 7695
rect 7380 7605 8100 7650
rect 8220 7620 8340 7650
rect 8700 7906 8820 7920
rect 7020 7320 7140 7334
rect 6870 7230 7140 7320
rect 6240 6990 6390 7080
rect 6810 7050 6900 7080
rect 6300 6810 6390 6990
rect 6600 6960 6900 7050
rect 7020 7095 7140 7110
rect 7020 7005 7740 7095
rect 7020 6990 7140 7005
rect 6300 6690 6420 6810
rect 6300 6480 6390 6690
rect 5580 6466 5820 6480
rect 5700 6390 5820 6466
rect 6240 6466 6480 6480
rect 5580 5280 5700 5294
rect 5820 6210 5970 6270
rect 5820 5340 5834 6210
rect 5956 5340 5970 6210
rect 5820 5190 5970 5340
rect 6240 5294 6300 6466
rect 6420 5294 6480 6466
rect 6870 6466 7140 6480
rect 6870 6390 7020 6466
rect 6240 5280 6480 5294
rect 6750 6210 6900 6270
rect 6750 5340 6764 6210
rect 6886 5340 6900 6210
rect 6750 5280 6900 5340
rect 7020 5280 7140 5294
rect 7980 5880 8100 7605
rect 8220 7290 8340 7410
rect 8700 7320 8820 7334
rect 8940 7906 9060 7920
rect 9180 7890 9300 8010
rect 9180 7440 9300 7470
rect 9420 7906 9540 7920
rect 9060 7334 9420 7350
rect 8940 7320 9540 7334
rect 9900 7906 10020 8010
rect 10290 7906 10410 7920
rect 9900 7320 10020 7334
rect 10140 7334 10290 7410
rect 10140 7320 10410 7334
rect 10860 7906 10980 7920
rect 10860 7320 10980 7334
rect 11100 7906 11220 7920
rect 11340 7890 11460 8010
rect 11340 7440 11460 7470
rect 11580 7906 11700 7920
rect 11220 7334 11580 7350
rect 11100 7320 11700 7334
rect 12300 7906 12420 8010
rect 12690 7906 12810 7920
rect 12300 7320 12420 7334
rect 12540 7334 12690 7410
rect 12540 7320 12810 7334
rect 13830 7906 13950 8010
rect 13830 7320 13950 7334
rect 14220 7906 14340 7920
rect 14460 7906 14580 8010
rect 14460 7620 14580 7634
rect 15420 7906 15540 8010
rect 15420 7620 15540 7634
rect 15660 7906 15780 7920
rect 15660 7620 15780 7634
rect 15900 7906 16020 8010
rect 15900 7620 16020 7634
rect 18060 7906 18180 8010
rect 18060 7620 18180 7634
rect 18300 7906 18420 7920
rect 18300 7620 18420 7634
rect 18540 7906 18660 8010
rect 18540 7620 18660 7634
rect 20700 7906 20820 8010
rect 14220 7320 14340 7334
rect 14460 7395 14580 7410
rect 8730 7110 8820 7320
rect 8970 7260 9510 7320
rect 8700 7095 9090 7110
rect 8580 7005 9090 7095
rect 9420 7095 9540 7110
rect 9420 7050 9900 7095
rect 9300 7020 9900 7050
rect 8700 6990 9090 7005
rect 9420 7005 9900 7020
rect 9420 6990 9540 7005
rect 8700 6495 8820 6510
rect 8340 6480 8820 6495
rect 9000 6480 9090 6990
rect 9180 6795 9300 6810
rect 9180 6705 9420 6795
rect 9180 6690 9300 6705
rect 8340 6405 8910 6480
rect 8700 6390 8910 6405
rect 9000 6466 9150 6480
rect 9000 6390 9030 6466
rect 8820 6210 8910 6390
rect 7980 5280 8100 5310
rect 6750 5190 6870 5280
rect 8220 5190 8340 5310
rect 8790 5866 8910 5880
rect 8790 5190 8910 5294
rect 9030 5280 9150 5294
rect 9420 6466 9540 6480
rect 9420 5190 9540 5294
rect 9900 5866 10020 5880
rect 9900 5190 10020 5294
rect 10140 5866 10260 7320
rect 10890 7110 10980 7320
rect 11130 7260 11670 7320
rect 10380 7095 10500 7110
rect 10860 7095 11250 7110
rect 10380 7005 11250 7095
rect 11580 7095 11700 7110
rect 12300 7095 12420 7110
rect 11580 7050 12420 7095
rect 11460 7020 12420 7050
rect 10380 6990 10500 7005
rect 10860 6990 11250 7005
rect 11580 7005 12420 7020
rect 11580 6990 11700 7005
rect 12300 6990 12420 7005
rect 10380 6390 10500 6510
rect 10860 6480 10980 6510
rect 11160 6480 11250 6990
rect 11340 6795 11460 6810
rect 11340 6705 12300 6795
rect 11340 6690 11460 6705
rect 11820 6495 11940 6510
rect 12540 6495 12660 7320
rect 13980 7095 14100 7110
rect 13140 7005 14100 7095
rect 13980 6990 14100 7005
rect 14220 6810 14310 7320
rect 14460 7305 15285 7395
rect 14460 7290 14580 7305
rect 15195 7095 15285 7305
rect 15690 7110 15780 7620
rect 16020 7305 16860 7395
rect 18060 7395 18180 7410
rect 16980 7305 18180 7395
rect 18060 7290 18180 7305
rect 18330 7110 18420 7620
rect 21090 7906 21210 7920
rect 20700 7320 20820 7334
rect 21060 7334 21090 7410
rect 21060 7320 21210 7334
rect 23340 7906 23460 8010
rect 26010 7920 26130 8010
rect 23730 7906 23850 7920
rect 23340 7320 23460 7334
rect 23580 7334 23730 7410
rect 25740 7906 25860 7920
rect 23850 7334 24300 7395
rect 15660 7095 15780 7110
rect 18300 7095 18420 7110
rect 15195 7005 15780 7095
rect 15660 6990 15780 7005
rect 13740 6795 13860 6810
rect 12900 6780 13860 6795
rect 14220 6795 14340 6810
rect 14460 6795 14580 6810
rect 12900 6750 13980 6780
rect 12900 6705 13860 6750
rect 13740 6690 13860 6705
rect 14220 6690 14580 6795
rect 10860 6390 11070 6480
rect 11160 6466 11310 6480
rect 11160 6390 11190 6466
rect 10980 6210 11070 6390
rect 10140 5280 10260 5294
rect 10380 5866 10500 5880
rect 10380 5190 10500 5294
rect 10950 5866 11070 5880
rect 10950 5190 11070 5294
rect 11190 5280 11310 5294
rect 11580 6466 11700 6480
rect 11820 6405 12660 6495
rect 11820 6390 11940 6405
rect 11580 5190 11700 5294
rect 12300 5866 12420 5880
rect 12300 5190 12420 5294
rect 12540 5866 12660 6405
rect 12780 6390 12900 6510
rect 14460 6480 14550 6690
rect 15690 6480 15780 6990
rect 17115 7005 18420 7095
rect 15900 6795 16020 6810
rect 17115 6795 17205 7005
rect 18300 6990 18420 7005
rect 18660 7005 20700 7095
rect 15900 6705 17205 6795
rect 15900 6690 16020 6705
rect 18330 6480 18420 6990
rect 13740 6466 14340 6480
rect 13740 6390 14220 6466
rect 13740 6346 13860 6390
rect 12540 5280 12660 5294
rect 12780 5866 12900 5880
rect 12780 5190 12900 5294
rect 13740 5280 13860 5324
rect 14220 5280 14340 5294
rect 14460 6466 14580 6480
rect 14460 5280 14580 5294
rect 15660 6360 15810 6480
rect 13980 5190 14100 5280
rect 15420 5190 15540 5310
rect 15810 5280 15930 5310
rect 18300 6360 18450 6480
rect 18060 5190 18180 5310
rect 18450 5280 18570 5310
rect 20700 5866 20820 5880
rect 20700 5190 20820 5294
rect 20940 5866 21060 7290
rect 23580 7305 24300 7334
rect 21300 7005 23340 7095
rect 21180 6495 21300 6510
rect 21180 6405 21420 6495
rect 21180 6390 21300 6405
rect 20940 5280 21060 5294
rect 21180 5866 21300 5880
rect 21180 5190 21300 5294
rect 23340 5866 23460 5880
rect 23340 5190 23460 5294
rect 23580 5866 23700 7305
rect 25980 7876 26130 7920
rect 25980 7454 25994 7876
rect 26116 7454 26130 7876
rect 25980 7410 26130 7454
rect 26400 7860 26640 7920
rect 26400 7440 26460 7860
rect 26580 7440 26640 7860
rect 26400 7380 26640 7440
rect 26910 7876 27060 8010
rect 26910 7454 26924 7876
rect 27046 7454 27060 7876
rect 26910 7410 27060 7454
rect 27180 7906 27300 7920
rect 25740 7320 25860 7334
rect 25740 7230 25950 7320
rect 26160 7170 26220 7260
rect 26160 7110 26250 7170
rect 25740 6990 25860 7110
rect 25980 7020 26250 7110
rect 26340 6870 26430 6960
rect 26160 6780 26430 6870
rect 26550 6870 26640 7380
rect 27180 7320 27300 7334
rect 27900 7906 28020 8010
rect 28290 7906 28410 7920
rect 27900 7320 28020 7334
rect 27060 7230 27300 7320
rect 28260 7334 28290 7410
rect 28260 7320 28410 7334
rect 29100 7906 29220 8010
rect 30330 7920 30450 8010
rect 29490 7906 29610 7920
rect 29100 7320 29220 7334
rect 29340 7334 29490 7410
rect 29340 7320 29610 7334
rect 30060 7906 30180 7920
rect 30300 7876 30450 7920
rect 30300 7454 30314 7876
rect 30436 7454 30450 7876
rect 30300 7410 30450 7454
rect 30720 7860 30960 7920
rect 30720 7440 30780 7860
rect 30900 7440 30960 7860
rect 30720 7380 30960 7440
rect 31230 7876 31380 8010
rect 31230 7454 31244 7876
rect 31366 7454 31380 7876
rect 31230 7410 31380 7454
rect 31500 7906 31620 7920
rect 30060 7320 30180 7334
rect 26760 7110 26850 7170
rect 27180 7095 27300 7110
rect 27180 7005 27660 7095
rect 27180 6990 27300 7005
rect 27900 6990 28020 7110
rect 26550 6810 26700 6870
rect 26550 6795 26820 6810
rect 26550 6780 27900 6795
rect 26610 6705 27900 6780
rect 26610 6690 26820 6705
rect 25980 6570 26370 6660
rect 23820 6495 23940 6510
rect 23820 6405 25260 6495
rect 23820 6390 23940 6405
rect 25980 6480 26070 6570
rect 26610 6480 26700 6690
rect 25740 6466 25950 6480
rect 23580 5280 23700 5294
rect 23820 5866 23940 5880
rect 23820 5190 23940 5294
rect 25860 6390 25950 6466
rect 26400 6466 26700 6480
rect 25740 5280 25860 5294
rect 25980 6210 26130 6270
rect 25980 5340 25994 6210
rect 26116 5340 26130 6210
rect 25980 5280 26130 5340
rect 26400 5294 26460 6466
rect 26580 6390 26700 6466
rect 26580 5294 26640 6390
rect 27060 6466 27300 6480
rect 27060 6390 27180 6466
rect 26400 5280 26640 5294
rect 26910 6210 27060 6270
rect 26910 5340 26924 6210
rect 27046 5340 27060 6210
rect 26010 5190 26130 5280
rect 26910 5190 27060 5340
rect 27180 5280 27300 5294
rect 27900 5866 28020 5880
rect 27900 5190 28020 5294
rect 28140 5866 28260 7290
rect 29100 7095 29220 7110
rect 28500 7005 29220 7095
rect 29100 6990 29220 7005
rect 29340 7095 29460 7320
rect 30060 7230 30330 7320
rect 30060 7095 30180 7110
rect 29340 7005 30180 7095
rect 28380 6390 28500 6510
rect 28140 5280 28260 5294
rect 28380 5866 28500 5880
rect 28380 5190 28500 5294
rect 29100 5866 29220 5880
rect 29100 5190 29220 5294
rect 29340 5866 29460 7005
rect 30060 6990 30180 7005
rect 30870 7080 30960 7380
rect 31500 7320 31620 7334
rect 31980 7906 32100 7920
rect 32220 7890 32340 8010
rect 32220 7440 32340 7470
rect 32460 7906 32580 7920
rect 32100 7334 32460 7350
rect 31980 7320 32580 7334
rect 32700 7906 32820 7920
rect 32700 7320 32820 7334
rect 33180 7906 33300 8010
rect 33570 7906 33690 7920
rect 33180 7320 33300 7334
rect 33420 7334 33570 7410
rect 33420 7320 33690 7334
rect 34710 7906 34830 7920
rect 35100 7906 35220 8010
rect 34830 7334 34980 7410
rect 34710 7320 34980 7334
rect 35100 7320 35220 7334
rect 36060 7906 36180 8010
rect 36450 7906 36570 7920
rect 36060 7320 36180 7334
rect 36300 7334 36450 7410
rect 37500 7906 37620 7920
rect 36900 7605 37500 7695
rect 37260 7395 37380 7410
rect 36570 7334 37380 7395
rect 31380 7230 31620 7320
rect 32010 7260 32550 7320
rect 30300 7050 30390 7080
rect 30300 6960 30600 7050
rect 30810 6990 30960 7080
rect 31080 7110 31170 7170
rect 31500 6990 31620 7110
rect 31740 7095 31860 7110
rect 31980 7095 32100 7110
rect 31740 7050 32100 7095
rect 32700 7110 32790 7320
rect 31740 7020 32220 7050
rect 31740 7005 32100 7020
rect 31740 6990 31860 7005
rect 31980 6990 32100 7005
rect 32430 6990 32460 7110
rect 32580 6990 32820 7110
rect 32940 7095 33060 7110
rect 33180 7095 33300 7110
rect 32940 7005 33300 7095
rect 32940 6990 33060 7005
rect 33180 6990 33300 7005
rect 30810 6810 30900 6990
rect 30780 6690 30900 6810
rect 31515 6795 31605 6990
rect 32220 6795 32340 6810
rect 31515 6705 32340 6795
rect 32220 6690 32340 6705
rect 30810 6480 30900 6690
rect 32430 6480 32520 6990
rect 33420 6795 33540 7320
rect 33420 6705 34005 6795
rect 32700 6495 32820 6510
rect 33180 6495 33300 6510
rect 32700 6480 33300 6495
rect 30060 6466 30330 6480
rect 29340 5280 29460 5294
rect 29580 5866 29700 5880
rect 29580 5190 29700 5294
rect 30180 6390 30330 6466
rect 30720 6466 30960 6480
rect 30060 5280 30180 5294
rect 30300 6210 30450 6270
rect 30300 5340 30314 6210
rect 30436 5340 30450 6210
rect 30300 5280 30450 5340
rect 30720 5294 30780 6466
rect 30900 5294 30960 6466
rect 31380 6466 31620 6480
rect 31380 6390 31500 6466
rect 30720 5280 30960 5294
rect 31230 6210 31380 6270
rect 31230 5340 31244 6210
rect 31366 5340 31380 6210
rect 30330 5190 30450 5280
rect 31230 5190 31380 5340
rect 31500 5280 31620 5294
rect 31980 6466 32100 6480
rect 31980 5190 32100 5294
rect 32370 6466 32520 6480
rect 32490 6390 32520 6466
rect 32610 6405 33300 6480
rect 32610 6390 32820 6405
rect 33180 6390 33300 6405
rect 32610 6210 32700 6390
rect 32370 5280 32490 5294
rect 32610 5866 32730 5880
rect 32610 5190 32730 5294
rect 33180 5866 33300 5880
rect 33180 5190 33300 5294
rect 33420 5866 33540 6705
rect 33915 6495 34005 6705
rect 34620 6495 34740 6510
rect 33915 6405 34740 6495
rect 34620 6390 34740 6405
rect 33420 5280 33540 5294
rect 33660 5866 33780 5880
rect 33660 5190 33780 5294
rect 34620 5866 34740 5880
rect 34620 5190 34740 5294
rect 34860 5866 34980 7320
rect 36300 7305 37380 7334
rect 37500 7320 37620 7334
rect 37740 7906 37860 7920
rect 37980 7890 38100 8010
rect 37980 7440 38100 7470
rect 38220 7906 38340 7920
rect 37860 7334 38220 7350
rect 37740 7320 38340 7334
rect 38940 7906 39060 8010
rect 39330 7906 39450 7920
rect 38940 7320 39060 7334
rect 39180 7334 39330 7410
rect 39180 7320 39450 7334
rect 40380 7906 40500 8010
rect 40770 7906 40890 7920
rect 40380 7320 40500 7334
rect 40620 7334 40770 7410
rect 43260 7906 43380 8010
rect 43260 7620 43380 7634
rect 43500 7906 43620 7920
rect 43500 7620 43620 7634
rect 43740 7906 43860 8010
rect 43740 7620 43860 7634
rect 44520 7906 44640 8010
rect 40620 7320 40890 7334
rect 36060 7095 36180 7110
rect 35460 7005 36180 7095
rect 36060 6990 36180 7005
rect 34860 5280 34980 5294
rect 35100 5866 35220 5880
rect 35100 5190 35220 5294
rect 36060 5866 36180 5880
rect 36060 5190 36180 5294
rect 36300 5866 36420 7305
rect 37260 7290 37380 7305
rect 37530 7110 37620 7320
rect 37770 7260 38310 7320
rect 37500 6990 37890 7110
rect 38220 7095 38340 7110
rect 38460 7095 38580 7110
rect 38220 7050 38580 7095
rect 38100 7020 38580 7050
rect 38220 7005 38580 7020
rect 38220 6990 38340 7005
rect 38460 6990 38580 7005
rect 38940 7095 39060 7110
rect 38820 7005 39060 7095
rect 38940 6990 39060 7005
rect 37500 6480 37620 6510
rect 37800 6480 37890 6990
rect 37980 6795 38100 6810
rect 38940 6795 39060 6810
rect 37980 6705 39060 6795
rect 37980 6690 38100 6705
rect 38940 6690 39060 6705
rect 38460 6495 38580 6510
rect 39180 6495 39300 7320
rect 39540 7005 39660 7095
rect 40380 7095 40500 7110
rect 39780 7005 40500 7095
rect 40380 6990 40500 7005
rect 37500 6390 37710 6480
rect 37800 6466 37950 6480
rect 37800 6390 37830 6466
rect 37620 6210 37710 6390
rect 36300 5280 36420 5294
rect 36540 5866 36660 5880
rect 36540 5190 36660 5294
rect 37590 5866 37710 5880
rect 37590 5190 37710 5294
rect 37830 5280 37950 5294
rect 38220 6466 38340 6480
rect 38460 6405 39300 6495
rect 38460 6390 38580 6405
rect 38220 5190 38340 5294
rect 38940 5866 39060 5880
rect 38940 5190 39060 5294
rect 39180 5866 39300 6405
rect 39420 6495 39540 6510
rect 40620 6495 40740 7320
rect 43260 7395 43380 7410
rect 42660 7305 43380 7395
rect 43260 7290 43380 7305
rect 43530 7110 43620 7620
rect 44520 7320 44640 7334
rect 44910 7906 45150 7920
rect 44910 7334 44970 7906
rect 45090 7334 45150 7906
rect 44910 7320 45150 7334
rect 45420 7906 45540 8010
rect 46620 7920 46740 8010
rect 45420 7320 45540 7334
rect 42180 7005 42540 7095
rect 43500 7095 43620 7110
rect 43500 7005 44220 7095
rect 43500 6990 43620 7005
rect 44700 6990 44820 7110
rect 39420 6405 40740 6495
rect 39420 6390 39540 6405
rect 39180 5280 39300 5294
rect 39420 5866 39540 5880
rect 39420 5190 39540 5294
rect 40380 5866 40500 5880
rect 40380 5190 40500 5294
rect 40620 5866 40740 6405
rect 43530 6480 43620 6990
rect 44970 6810 45060 7320
rect 45180 7095 45300 7110
rect 46380 7095 46500 7650
rect 46620 7620 46740 7650
rect 47340 7906 47460 7920
rect 46620 7290 46740 7410
rect 47340 7320 47460 7334
rect 47580 7906 47700 7920
rect 47820 7890 47940 8010
rect 47820 7440 47940 7470
rect 48060 7906 48180 7920
rect 47700 7334 48060 7350
rect 47580 7320 48180 7334
rect 47370 7110 47460 7320
rect 47610 7260 48150 7320
rect 45180 7005 46500 7095
rect 45180 6990 45300 7005
rect 45180 6930 45270 6990
rect 43740 6795 43860 6810
rect 43740 6705 43980 6795
rect 43740 6690 43860 6705
rect 44580 6750 44700 6780
rect 44940 6690 45060 6810
rect 44970 6660 45060 6690
rect 45420 6690 45540 6810
rect 44970 6570 45270 6660
rect 45180 6480 45270 6570
rect 40620 5280 40740 5294
rect 40860 5866 40980 5880
rect 40860 5190 40980 5294
rect 43500 6360 43650 6480
rect 43260 5190 43380 5310
rect 43650 5280 43770 5310
rect 44460 6466 45060 6480
rect 44460 6390 44940 6466
rect 44460 6346 44580 6390
rect 44460 5280 44580 5324
rect 45420 6466 45540 6480
rect 45060 5294 45420 5370
rect 44940 5280 45540 5294
rect 46380 5880 46500 7005
rect 46620 7095 46740 7110
rect 47340 7095 47730 7110
rect 46620 7005 47730 7095
rect 47940 7020 48060 7050
rect 46620 6990 46740 7005
rect 47340 6990 47730 7005
rect 47640 6480 47730 6990
rect 47460 6210 47550 6480
rect 47640 6466 47790 6480
rect 47640 6390 47670 6466
rect 46380 5280 46500 5310
rect 44700 5190 44820 5280
rect 46620 5190 46740 5310
rect 47430 5866 47550 5880
rect 47430 5190 47550 5294
rect 47670 5280 47790 5294
rect 48060 6466 48180 6480
rect 48060 5190 48180 5294
rect 1155 5160 54240 5190
rect 1155 5040 1214 5160
rect 2086 5040 5220 5160
rect 5340 5040 5460 5160
rect 5580 5040 5700 5160
rect 5820 5040 6180 5160
rect 6300 5040 6660 5160
rect 6780 5040 7140 5160
rect 7260 5040 7380 5160
rect 7500 5040 7620 5160
rect 7740 5040 7860 5160
rect 7980 5040 8340 5160
rect 8460 5040 8580 5160
rect 8700 5040 9060 5160
rect 9180 5040 9540 5160
rect 9660 5040 9780 5160
rect 9900 5040 10260 5160
rect 10380 5040 10500 5160
rect 10620 5040 10740 5160
rect 10860 5040 11220 5160
rect 11340 5040 11700 5160
rect 11820 5040 11940 5160
rect 12060 5040 12180 5160
rect 12300 5040 12660 5160
rect 12780 5040 12900 5160
rect 13020 5040 13140 5160
rect 13260 5040 13380 5160
rect 13500 5040 13620 5160
rect 13740 5040 14100 5160
rect 14220 5040 14580 5160
rect 14700 5040 14820 5160
rect 14940 5040 15060 5160
rect 15180 5040 15300 5160
rect 15420 5040 15780 5160
rect 15900 5040 16020 5160
rect 16140 5040 16260 5160
rect 16380 5040 16500 5160
rect 16620 5040 16740 5160
rect 16860 5040 16980 5160
rect 17100 5040 17220 5160
rect 17340 5040 17460 5160
rect 17580 5040 17700 5160
rect 17820 5040 17940 5160
rect 18060 5040 18420 5160
rect 18540 5040 18660 5160
rect 18780 5040 18900 5160
rect 19020 5040 19140 5160
rect 19260 5040 19380 5160
rect 19500 5040 19620 5160
rect 19740 5040 19860 5160
rect 19980 5040 20100 5160
rect 20220 5040 20340 5160
rect 20460 5040 20580 5160
rect 20700 5040 21060 5160
rect 21180 5040 21300 5160
rect 21420 5040 21540 5160
rect 21660 5040 21780 5160
rect 21900 5040 22020 5160
rect 22140 5040 22260 5160
rect 22380 5040 22500 5160
rect 22620 5040 22740 5160
rect 22860 5040 22980 5160
rect 23100 5040 23220 5160
rect 23340 5040 23700 5160
rect 23820 5040 23940 5160
rect 24060 5040 24180 5160
rect 24300 5040 24420 5160
rect 24540 5040 24660 5160
rect 24780 5040 24900 5160
rect 25020 5040 25140 5160
rect 25260 5040 25380 5160
rect 25500 5040 25620 5160
rect 25740 5040 26100 5160
rect 26220 5040 26580 5160
rect 26700 5040 27060 5160
rect 27180 5040 27300 5160
rect 27420 5040 27540 5160
rect 27660 5040 27780 5160
rect 27900 5040 28260 5160
rect 28380 5040 28500 5160
rect 28620 5040 28740 5160
rect 28860 5040 28980 5160
rect 29100 5040 29460 5160
rect 29580 5040 29700 5160
rect 29820 5040 29940 5160
rect 30060 5040 30420 5160
rect 30540 5040 30900 5160
rect 31020 5040 31380 5160
rect 31500 5040 31620 5160
rect 31740 5040 31860 5160
rect 31980 5040 32340 5160
rect 32460 5040 32820 5160
rect 32940 5040 33060 5160
rect 33180 5040 33540 5160
rect 33660 5040 33780 5160
rect 33900 5040 34020 5160
rect 34140 5040 34260 5160
rect 34380 5040 34500 5160
rect 34620 5040 34740 5160
rect 34860 5040 35220 5160
rect 35340 5040 35460 5160
rect 35580 5040 35700 5160
rect 35820 5040 35940 5160
rect 36060 5040 36420 5160
rect 36540 5040 36660 5160
rect 36780 5040 36900 5160
rect 37020 5040 37140 5160
rect 37260 5040 37380 5160
rect 37500 5040 37860 5160
rect 37980 5040 38340 5160
rect 38460 5040 38580 5160
rect 38700 5040 38820 5160
rect 38940 5040 39300 5160
rect 39420 5040 39540 5160
rect 39660 5040 39780 5160
rect 39900 5040 40020 5160
rect 40140 5040 40260 5160
rect 40380 5040 40740 5160
rect 40860 5040 40980 5160
rect 41100 5040 41220 5160
rect 41340 5040 41460 5160
rect 41580 5040 41700 5160
rect 41820 5040 41940 5160
rect 42060 5040 42180 5160
rect 42300 5040 42420 5160
rect 42540 5040 42660 5160
rect 42780 5040 42900 5160
rect 43020 5040 43140 5160
rect 43260 5040 43620 5160
rect 43740 5040 43860 5160
rect 43980 5040 44100 5160
rect 44220 5040 44340 5160
rect 44460 5040 44820 5160
rect 44940 5040 45300 5160
rect 45420 5040 45540 5160
rect 45660 5040 45780 5160
rect 45900 5040 46020 5160
rect 46140 5040 46260 5160
rect 46380 5040 46740 5160
rect 46860 5040 46980 5160
rect 47100 5040 47220 5160
rect 47340 5040 47700 5160
rect 47820 5040 48180 5160
rect 48300 5040 48420 5160
rect 48540 5040 48660 5160
rect 48780 5040 48900 5160
rect 49020 5040 49140 5160
rect 49260 5040 49380 5160
rect 49500 5040 49620 5160
rect 49740 5040 49860 5160
rect 49980 5040 50100 5160
rect 50220 5040 53310 5160
rect 54180 5040 54240 5160
rect 1155 5010 54240 5040
rect 3135 3976 52260 4035
rect 3135 3104 3194 3976
rect 4066 3104 51330 3976
rect 52200 3104 52260 3976
rect 3135 3045 52260 3104
rect 17220 2805 35580 2895
rect 17460 2505 28620 2595
rect 18660 2205 21180 2295
rect 1155 1996 54240 2055
rect 1155 1124 1214 1996
rect 2086 1124 53310 1996
rect 54180 1124 54240 1996
rect 1155 1065 54240 1124
<< m2contact >>
rect 1214 47204 2086 48076
rect 53310 47204 54180 48076
rect 15300 46590 15420 46710
rect 32940 46590 33060 46710
rect 3194 45224 4066 46096
rect 51330 45224 52200 46096
rect 3194 44040 4066 44160
rect 51330 44040 52200 44160
rect 5340 42990 5460 43110
rect 9210 43200 9330 43320
rect 9420 43170 9540 43290
rect 8940 42990 9060 43110
rect 9930 43170 10050 43290
rect 10140 43200 10260 43320
rect 7260 42390 7380 42510
rect 12780 43290 12900 43410
rect 10620 42990 10740 43110
rect 12780 42990 12900 43110
rect 14220 42990 14340 43110
rect 8700 42690 8820 42810
rect 9390 42660 9510 42780
rect 10860 42690 10980 42810
rect 11580 42690 11700 42810
rect 13020 42690 13140 42810
rect 17100 42990 17220 43110
rect 19500 43200 19620 43320
rect 19710 43170 19830 43290
rect 17580 42990 17700 43110
rect 19260 42990 19380 43110
rect 9210 42360 9330 42480
rect 10140 42360 10260 42480
rect 20220 43170 20340 43290
rect 20490 43200 20610 43320
rect 20940 43290 21060 43410
rect 20100 42960 20220 43080
rect 18060 42690 18180 42810
rect 22890 43200 23010 43320
rect 23100 43170 23220 43290
rect 22620 42990 22740 43110
rect 31500 43590 31620 43710
rect 23610 43170 23730 43290
rect 23820 43200 23940 43320
rect 25740 42990 25860 43110
rect 18780 42390 18900 42510
rect 19500 42360 19620 42480
rect 20490 42360 20610 42480
rect 23070 42660 23190 42780
rect 26220 42690 26340 42810
rect 27180 42990 27300 43110
rect 27900 42990 28020 43110
rect 28140 42690 28260 42810
rect 22890 42360 23010 42480
rect 23820 42360 23940 42480
rect 27180 42390 27300 42510
rect 29580 42990 29700 43110
rect 31260 42990 31380 43110
rect 34620 43290 34740 43410
rect 36090 43200 36210 43320
rect 36300 43170 36420 43290
rect 33660 42990 33780 43110
rect 35820 42990 35940 43110
rect 36810 43170 36930 43290
rect 37020 43200 37140 43320
rect 33180 42390 33300 42510
rect 39660 43200 39780 43320
rect 39870 43170 39990 43290
rect 39420 42990 39540 43110
rect 40380 43170 40500 43290
rect 40590 43200 40710 43320
rect 35340 42690 35460 42810
rect 36270 42660 36390 42780
rect 36090 42360 36210 42480
rect 37020 42360 37140 42480
rect 37740 42390 37860 42510
rect 38220 42690 38340 42810
rect 40860 42990 40980 43110
rect 40410 42660 40530 42780
rect 42300 42990 42420 43110
rect 44940 42990 45060 43110
rect 39660 42360 39780 42480
rect 40590 42360 40710 42480
rect 43980 42390 44100 42510
rect 45420 43290 45540 43410
rect 45930 43200 46050 43320
rect 46140 43170 46260 43290
rect 46650 43170 46770 43290
rect 46860 43200 46980 43320
rect 47610 43200 47730 43320
rect 47820 43170 47940 43290
rect 47100 42990 47220 43110
rect 47340 42990 47460 43110
rect 48330 43170 48450 43290
rect 48540 43200 48660 43320
rect 48780 42990 48900 43110
rect 44940 42390 45060 42510
rect 46110 42660 46230 42780
rect 47790 42660 47910 42780
rect 54434 42690 54556 42810
rect 45930 42360 46050 42480
rect 46860 42360 46980 42480
rect 47610 42360 47730 42480
rect 48540 42360 48660 42480
rect 1214 41040 2086 41160
rect 53310 41040 54180 41160
rect 7260 40590 7380 40710
rect 5580 39390 5700 39510
rect 7020 38790 7140 38910
rect 10140 39690 10260 39810
rect 11790 39720 11910 39840
rect 12780 39720 12900 39840
rect 9660 39090 9780 39210
rect 10380 38790 10500 38910
rect 11340 39390 11460 39510
rect 13980 39690 14100 39810
rect 11580 39090 11700 39210
rect 12180 39120 12300 39240
rect 11790 38880 11910 39000
rect 12060 38910 12180 39030
rect 13500 39090 13620 39210
rect 12570 38910 12690 39030
rect 12780 38880 12900 39000
rect 15660 39690 15780 39810
rect 15180 39090 15300 39210
rect 15420 38790 15540 38910
rect 17340 39690 17460 39810
rect 17580 39690 17700 39810
rect 16140 39090 16260 39210
rect 18780 39390 18900 39510
rect 20940 39690 21060 39810
rect 22170 39720 22290 39840
rect 23100 39720 23220 39840
rect 19740 39090 19860 39210
rect 19020 38790 19140 38910
rect 22350 39420 22470 39540
rect 21420 39090 21540 39210
rect 21660 39090 21780 39210
rect 21900 39090 22020 39210
rect 24300 39390 24420 39510
rect 25740 39690 25860 39810
rect 26220 39390 26340 39510
rect 22170 38880 22290 39000
rect 22380 38910 22500 39030
rect 24060 39090 24180 39210
rect 24780 39090 24900 39210
rect 22890 38910 23010 39030
rect 23100 38880 23220 39000
rect 29580 39690 29700 39810
rect 31260 39090 31380 39210
rect 33690 39720 33810 39840
rect 34620 39720 34740 39840
rect 33870 39420 33990 39540
rect 35340 39390 35460 39510
rect 32460 39090 32580 39210
rect 33690 38880 33810 39000
rect 33900 38910 34020 39030
rect 34860 39090 34980 39210
rect 37260 39690 37380 39810
rect 34410 38910 34530 39030
rect 34620 38880 34740 39000
rect 38700 39390 38820 39510
rect 38220 39090 38340 39210
rect 39420 39090 39540 39210
rect 40860 39690 40980 39810
rect 41580 38790 41700 38910
rect 43740 39690 43860 39810
rect 45180 39690 45300 39810
rect 42540 39090 42660 39210
rect 43980 39090 44100 39210
rect 44700 38790 44820 38910
rect 46620 39390 46740 39510
rect 47820 39390 47940 39510
rect 46140 39090 46260 39210
rect 46860 39090 46980 39210
rect 49740 39090 49860 39210
rect 3194 38040 4066 38160
rect 51330 38040 52200 38160
rect 7020 37590 7140 37710
rect 7500 37590 7620 37710
rect 7500 37290 7620 37410
rect 13500 37590 13620 37710
rect 8460 36990 8580 37110
rect 15900 36990 16020 37110
rect 11340 36390 11460 36510
rect 11820 36390 11940 36510
rect 12060 36390 12180 36510
rect 13740 36690 13860 36810
rect 13020 36390 13140 36510
rect 15660 36690 15780 36810
rect 17340 36990 17460 37110
rect 17580 36990 17700 37110
rect 17100 36390 17220 36510
rect 17820 36390 17940 36510
rect 19500 36990 19620 37110
rect 18540 36390 18660 36510
rect 21180 37290 21300 37410
rect 22380 36990 22500 37110
rect 23820 37290 23940 37410
rect 22860 36390 22980 36510
rect 25020 36390 25140 36510
rect 25500 36990 25620 37110
rect 27420 36990 27540 37110
rect 25500 36690 25620 36810
rect 27180 36690 27300 36810
rect 29100 36990 29220 37110
rect 28860 36390 28980 36510
rect 30060 36990 30180 37110
rect 30300 36690 30420 36810
rect 29580 36390 29700 36510
rect 32940 37290 33060 37410
rect 31740 36990 31860 37110
rect 32700 36990 32820 37110
rect 31980 36390 32100 36510
rect 34860 37290 34980 37410
rect 34380 36990 34500 37110
rect 34620 36990 34740 37110
rect 35820 37200 35940 37320
rect 36030 37170 36150 37290
rect 36540 37170 36660 37290
rect 36750 37200 36870 37320
rect 37260 37290 37380 37410
rect 37020 36990 37140 37110
rect 40350 37590 40470 37710
rect 35100 36390 35220 36510
rect 36570 36660 36690 36780
rect 35820 36360 35940 36480
rect 36750 36360 36870 36480
rect 41100 37290 41220 37410
rect 40620 36990 40740 37110
rect 39420 36690 39540 36810
rect 40860 36690 40980 36810
rect 42060 36990 42180 37110
rect 42300 36390 42420 36510
rect 43740 37290 43860 37410
rect 43980 36990 44100 37110
rect 44700 36690 44820 36810
rect 47580 36990 47700 37110
rect 46620 36390 46740 36510
rect 49740 36990 49860 37110
rect 1214 35040 2086 35160
rect 53310 35040 54180 35160
rect 5820 33690 5940 33810
rect 9150 33720 9270 33840
rect 10140 33720 10260 33840
rect 11310 33720 11430 33840
rect 12300 33720 12420 33840
rect 7020 33390 7140 33510
rect 8220 33390 8340 33510
rect 6540 33090 6660 33210
rect 7260 33090 7380 33210
rect 7500 33090 7620 33210
rect 8700 33090 8820 33210
rect 9540 33120 9660 33240
rect 9150 32880 9270 33000
rect 9420 32910 9540 33030
rect 10860 33090 10980 33210
rect 11700 33120 11820 33240
rect 9930 32910 10050 33030
rect 10140 32880 10260 33000
rect 11310 32880 11430 33000
rect 11580 32910 11700 33030
rect 12090 32910 12210 33030
rect 12300 32880 12420 33000
rect 13980 33990 14100 34110
rect 13980 32790 14100 32910
rect 14940 32790 15060 32910
rect 15660 33690 15780 33810
rect 18300 33690 18420 33810
rect 16380 33090 16500 33210
rect 19980 33090 20100 33210
rect 22860 33390 22980 33510
rect 23340 33390 23460 33510
rect 23580 33390 23700 33510
rect 24060 33390 24180 33510
rect 25500 33690 25620 33810
rect 26250 33720 26370 33840
rect 27180 33720 27300 33840
rect 26430 33420 26550 33540
rect 22620 33090 22740 33210
rect 24300 33090 24420 33210
rect 25260 33090 25380 33210
rect 26250 32880 26370 33000
rect 26460 32910 26580 33030
rect 27420 33090 27540 33210
rect 26970 32910 27090 33030
rect 27180 32880 27300 33000
rect 31020 33690 31140 33810
rect 30540 32790 30660 32910
rect 31500 33390 31620 33510
rect 31980 33390 32100 33510
rect 31500 33090 31620 33210
rect 31740 33090 31860 33210
rect 32940 33090 33060 33210
rect 34620 33090 34740 33210
rect 35100 33690 35220 33810
rect 35340 33090 35460 33210
rect 38700 33990 38820 34110
rect 37980 33090 38100 33210
rect 38220 33090 38340 33210
rect 39420 33690 39540 33810
rect 40380 33390 40500 33510
rect 41580 33690 41700 33810
rect 41340 33090 41460 33210
rect 42060 33690 42180 33810
rect 44490 33720 44610 33840
rect 45420 33720 45540 33840
rect 44670 33420 44790 33540
rect 45900 33390 46020 33510
rect 43500 33090 43620 33210
rect 47580 33690 47700 33810
rect 44490 32880 44610 33000
rect 44700 32910 44820 33030
rect 45660 33090 45780 33210
rect 46140 33090 46260 33210
rect 45210 32910 45330 33030
rect 45420 32880 45540 33000
rect 48060 33390 48180 33510
rect 48060 33090 48180 33210
rect 48300 33090 48420 33210
rect 49500 33090 49620 33210
rect 3194 32040 4066 32160
rect 51330 32040 52200 32160
rect 5580 31200 5700 31320
rect 5790 31170 5910 31290
rect 5340 30990 5460 31110
rect 6300 31170 6420 31290
rect 6570 31200 6690 31320
rect 6180 30960 6300 31080
rect 7020 30990 7140 31110
rect 8460 30990 8580 31110
rect 5580 30360 5700 30480
rect 6570 30360 6690 30480
rect 8940 30390 9060 30510
rect 9180 30390 9300 30510
rect 11370 31200 11490 31320
rect 11580 31170 11700 31290
rect 10140 30990 10260 31110
rect 11100 30990 11220 31110
rect 12090 31170 12210 31290
rect 12300 31200 12420 31320
rect 14910 31200 15030 31320
rect 15180 31170 15300 31290
rect 12780 30990 12900 31110
rect 13980 30990 14100 31110
rect 15300 30960 15420 31080
rect 11550 30660 11670 30780
rect 15690 31170 15810 31290
rect 15900 31200 16020 31320
rect 17310 31200 17430 31320
rect 17580 31170 17700 31290
rect 16860 30990 16980 31110
rect 17100 30990 17220 31110
rect 17700 30960 17820 31080
rect 18090 31170 18210 31290
rect 18300 31200 18420 31320
rect 19530 31200 19650 31320
rect 19740 31170 19860 31290
rect 19020 30990 19140 31110
rect 19260 30990 19380 31110
rect 23580 31590 23700 31710
rect 20250 31170 20370 31290
rect 20460 31200 20580 31320
rect 21180 30990 21300 31110
rect 19710 30660 19830 30780
rect 11370 30360 11490 30480
rect 12300 30360 12420 30480
rect 14910 30360 15030 30480
rect 15900 30360 16020 30480
rect 17310 30360 17430 30480
rect 18300 30360 18420 30480
rect 19530 30360 19650 30480
rect 20460 30360 20580 30480
rect 22140 30990 22260 31110
rect 22860 30990 22980 31110
rect 21660 30390 21780 30510
rect 22620 30690 22740 30810
rect 24300 31290 24420 31410
rect 25740 31590 25860 31710
rect 24060 30090 24180 30210
rect 25740 30990 25860 31110
rect 26700 30990 26820 31110
rect 25260 30390 25380 30510
rect 25740 30390 25860 30510
rect 25980 30390 26100 30510
rect 28620 31290 28740 31410
rect 28380 30990 28500 31110
rect 31020 31200 31140 31320
rect 31230 31170 31350 31290
rect 29820 30990 29940 31110
rect 30060 30990 30180 31110
rect 31740 31170 31860 31290
rect 31950 31200 32070 31320
rect 33420 31290 33540 31410
rect 29100 30390 29220 30510
rect 32220 30990 32340 31110
rect 33180 30990 33300 31110
rect 31770 30660 31890 30780
rect 31020 30360 31140 30480
rect 31950 30360 32070 30480
rect 33900 30990 34020 31110
rect 35820 31290 35940 31410
rect 35100 30990 35220 31110
rect 36540 30690 36660 30810
rect 37500 30090 37620 30210
rect 38460 30990 38580 31110
rect 38220 30390 38340 30510
rect 41340 31290 41460 31410
rect 45660 31590 45780 31710
rect 40860 30390 40980 30510
rect 41580 30390 41700 30510
rect 43260 30990 43380 31110
rect 43740 30990 43860 31110
rect 43980 30990 44100 31110
rect 43500 30690 43620 30810
rect 43980 30690 44100 30810
rect 48330 31200 48450 31320
rect 48540 31170 48660 31290
rect 46620 30990 46740 31110
rect 47340 30990 47460 31110
rect 49050 31170 49170 31290
rect 49260 31200 49380 31320
rect 49740 30990 49860 31110
rect 46140 30390 46260 30510
rect 48510 30660 48630 30780
rect 49500 30690 49620 30810
rect 48330 30360 48450 30480
rect 49260 30360 49380 30480
rect 1214 29040 2086 29160
rect 53310 29040 54180 29160
rect 7290 27720 7410 27840
rect 8220 27720 8340 27840
rect 7470 27420 7590 27540
rect 7020 27090 7140 27210
rect 7290 26880 7410 27000
rect 7500 26910 7620 27030
rect 8460 27090 8580 27210
rect 8700 27090 8820 27210
rect 8010 26910 8130 27030
rect 8220 26880 8340 27000
rect 9180 27690 9300 27810
rect 9660 27720 9780 27840
rect 10650 27720 10770 27840
rect 9180 27090 9300 27210
rect 9660 26880 9780 27000
rect 9870 26910 9990 27030
rect 11340 27390 11460 27510
rect 10260 27120 10380 27240
rect 11820 27090 11940 27210
rect 12060 27090 12180 27210
rect 10380 26910 10500 27030
rect 10650 26880 10770 27000
rect 14460 27990 14580 28110
rect 15180 27090 15300 27210
rect 15420 27090 15540 27210
rect 16380 27690 16500 27810
rect 16620 27690 16740 27810
rect 17820 27090 17940 27210
rect 18780 27690 18900 27810
rect 19260 27690 19380 27810
rect 19740 27390 19860 27510
rect 18300 26790 18420 26910
rect 20940 27090 21060 27210
rect 21420 27690 21540 27810
rect 21660 27090 21780 27210
rect 22860 27990 22980 28110
rect 23580 27690 23700 27810
rect 23100 27090 23220 27210
rect 23580 27090 23700 27210
rect 24060 27090 24180 27210
rect 25500 27690 25620 27810
rect 27180 27690 27300 27810
rect 27900 27690 28020 27810
rect 25500 27090 25620 27210
rect 29340 27690 29460 27810
rect 30300 27690 30420 27810
rect 33210 27720 33330 27840
rect 34140 27720 34260 27840
rect 28620 27090 28740 27210
rect 29100 27090 29220 27210
rect 33390 27420 33510 27540
rect 30780 27090 30900 27210
rect 32460 27090 32580 27210
rect 32700 27090 32820 27210
rect 33210 26880 33330 27000
rect 33420 26910 33540 27030
rect 18780 26490 18900 26610
rect 34620 27090 34740 27210
rect 33930 26910 34050 27030
rect 34140 26880 34260 27000
rect 35340 27690 35460 27810
rect 35580 27090 35700 27210
rect 37020 27690 37140 27810
rect 37260 27690 37380 27810
rect 37500 27690 37620 27810
rect 38700 27090 38820 27210
rect 39420 27690 39540 27810
rect 39930 27720 40050 27840
rect 40860 27720 40980 27840
rect 40110 27420 40230 27540
rect 39180 27090 39300 27210
rect 42060 27690 42180 27810
rect 39930 26880 40050 27000
rect 40140 26910 40260 27030
rect 41100 27090 41220 27210
rect 40650 26910 40770 27030
rect 40860 26880 40980 27000
rect 43500 27390 43620 27510
rect 44700 27390 44820 27510
rect 45180 27690 45300 27810
rect 46140 27390 46260 27510
rect 42780 27090 42900 27210
rect 43740 27090 43860 27210
rect 44460 27090 44580 27210
rect 44940 27090 45060 27210
rect 45900 27090 46020 27210
rect 47340 27390 47460 27510
rect 48540 27090 48660 27210
rect 49020 27690 49140 27810
rect 49020 27090 49140 27210
rect 49260 27090 49380 27210
rect 49740 27090 49860 27210
rect 3194 26040 4066 26160
rect 51330 26040 52200 26160
rect 5610 25200 5730 25320
rect 5820 25170 5940 25290
rect 6330 25170 6450 25290
rect 6540 25200 6660 25320
rect 6780 24990 6900 25110
rect 5790 24660 5910 24780
rect 8460 24990 8580 25110
rect 5610 24360 5730 24480
rect 6540 24360 6660 24480
rect 9690 25200 9810 25320
rect 9900 25170 10020 25290
rect 9180 24990 9300 25110
rect 9420 24990 9540 25110
rect 10410 25170 10530 25290
rect 10620 25200 10740 25320
rect 9870 24660 9990 24780
rect 9180 24390 9300 24510
rect 9690 24360 9810 24480
rect 10620 24360 10740 24480
rect 15660 24990 15780 25110
rect 13980 24390 14100 24510
rect 15420 24690 15540 24810
rect 18780 24390 18900 24510
rect 19740 24390 19860 24510
rect 23340 25290 23460 25410
rect 21180 24990 21300 25110
rect 21900 24990 22020 25110
rect 25740 25200 25860 25320
rect 25950 25170 26070 25290
rect 26460 25170 26580 25290
rect 26670 25200 26790 25320
rect 27420 24990 27540 25110
rect 29340 24990 29460 25110
rect 23580 24690 23700 24810
rect 24540 24690 24660 24810
rect 26490 24660 26610 24780
rect 25740 24360 25860 24480
rect 26670 24360 26790 24480
rect 27900 24390 28020 24510
rect 31740 24990 31860 25110
rect 30780 24390 30900 24510
rect 31020 24390 31140 24510
rect 32460 25290 32580 25410
rect 32460 24690 32580 24810
rect 34620 24990 34740 25110
rect 34620 24390 34740 24510
rect 35820 25290 35940 25410
rect 36060 24990 36180 25110
rect 35100 24390 35220 24510
rect 36540 24990 36660 25110
rect 36540 24390 36660 24510
rect 36780 24390 36900 24510
rect 39420 24390 39540 24510
rect 42540 25290 42660 25410
rect 44700 25590 44820 25710
rect 43980 25290 44100 25410
rect 42300 24390 42420 24510
rect 43740 24690 43860 24810
rect 48090 25200 48210 25320
rect 48300 25170 48420 25290
rect 47820 24990 47940 25110
rect 48810 25170 48930 25290
rect 49020 25200 49140 25320
rect 49500 24990 49620 25110
rect 48270 24660 48390 24780
rect 48090 24360 48210 24480
rect 49020 24360 49140 24480
rect 1214 23040 2086 23160
rect 53310 23040 54180 23160
rect 5610 21720 5730 21840
rect 6540 21720 6660 21840
rect 5790 21420 5910 21540
rect 5610 20880 5730 21000
rect 5820 20910 5940 21030
rect 6780 21090 6900 21210
rect 6330 20910 6450 21030
rect 6540 20880 6660 21000
rect 9660 21390 9780 21510
rect 8940 21090 9060 21210
rect 10140 21690 10260 21810
rect 14490 21720 14610 21840
rect 15420 21720 15540 21840
rect 11580 21390 11700 21510
rect 14670 21420 14790 21540
rect 10380 21090 10500 21210
rect 12300 21090 12420 21210
rect 14220 21090 14340 21210
rect 14490 20880 14610 21000
rect 14700 20910 14820 21030
rect 15660 21090 15780 21210
rect 15210 20910 15330 21030
rect 15420 20880 15540 21000
rect 18060 21090 18180 21210
rect 18540 21690 18660 21810
rect 19020 21720 19140 21840
rect 19950 21720 20070 21840
rect 20700 21720 20820 21840
rect 21630 21720 21750 21840
rect 19770 21420 19890 21540
rect 22140 21690 22260 21810
rect 21450 21420 21570 21540
rect 18780 21090 18900 21210
rect 17820 20790 17940 20910
rect 16860 20490 16980 20610
rect 18300 20790 18420 20910
rect 19020 20880 19140 21000
rect 19230 20910 19350 21030
rect 20220 21090 20340 21210
rect 20460 21090 20580 21210
rect 22620 21390 22740 21510
rect 25980 21690 26100 21810
rect 19740 20910 19860 21030
rect 19950 20880 20070 21000
rect 20700 20880 20820 21000
rect 20910 20910 21030 21030
rect 21900 21090 22020 21210
rect 22380 21090 22500 21210
rect 21420 20910 21540 21030
rect 21630 20880 21750 21000
rect 24300 20790 24420 20910
rect 28380 21390 28500 21510
rect 27420 21090 27540 21210
rect 28140 21090 28260 21210
rect 29820 21690 29940 21810
rect 29580 21390 29700 21510
rect 30780 21090 30900 21210
rect 31260 21090 31380 21210
rect 32460 21690 32580 21810
rect 32940 21090 33060 21210
rect 33660 21690 33780 21810
rect 34620 21090 34740 21210
rect 33420 20790 33540 20910
rect 35100 21690 35220 21810
rect 36540 21690 36660 21810
rect 37050 21720 37170 21840
rect 37980 21720 38100 21840
rect 35340 21090 35460 21210
rect 34860 20790 34980 20910
rect 37230 21420 37350 21540
rect 37050 20880 37170 21000
rect 37260 20910 37380 21030
rect 37770 20910 37890 21030
rect 37980 20880 38100 21000
rect 39660 21090 39780 21210
rect 40380 21090 40500 21210
rect 41100 21690 41220 21810
rect 44490 21720 44610 21840
rect 45420 21720 45540 21840
rect 46140 21720 46260 21840
rect 47070 21720 47190 21840
rect 44670 21420 44790 21540
rect 42300 21090 42420 21210
rect 43500 21090 43620 21210
rect 43740 21090 43860 21210
rect 46890 21420 47010 21540
rect 44490 20880 44610 21000
rect 44700 20910 44820 21030
rect 45900 21090 46020 21210
rect 45210 20910 45330 21030
rect 45420 20880 45540 21000
rect 46140 20880 46260 21000
rect 46350 20910 46470 21030
rect 47340 21090 47460 21210
rect 49980 21390 50100 21510
rect 46860 20910 46980 21030
rect 47070 20880 47190 21000
rect 47580 20790 47700 20910
rect 49740 21090 49860 21210
rect 3194 20040 4066 20160
rect 51330 20040 52200 20160
rect 5340 19590 5460 19710
rect 9180 19200 9300 19320
rect 9390 19170 9510 19290
rect 6780 18990 6900 19110
rect 8940 18990 9060 19110
rect 9900 19170 10020 19290
rect 10110 19200 10230 19320
rect 11790 19200 11910 19320
rect 12060 19170 12180 19290
rect 5580 18390 5700 18510
rect 6060 18690 6180 18810
rect 10380 18990 10500 19110
rect 11100 18990 11220 19110
rect 12180 18960 12300 19080
rect 9930 18660 10050 18780
rect 12570 19170 12690 19290
rect 12780 19200 12900 19320
rect 13770 19200 13890 19320
rect 13980 19170 14100 19290
rect 13260 18990 13380 19110
rect 13500 18990 13620 19110
rect 14490 19170 14610 19290
rect 14700 19200 14820 19320
rect 15660 18990 15780 19110
rect 13950 18660 14070 18780
rect 16860 19290 16980 19410
rect 19740 19290 19860 19410
rect 19500 18990 19620 19110
rect 9180 18360 9300 18480
rect 10110 18360 10230 18480
rect 11790 18360 11910 18480
rect 12780 18360 12900 18480
rect 13770 18360 13890 18480
rect 14700 18360 14820 18480
rect 16380 18390 16500 18510
rect 20940 18990 21060 19110
rect 20220 18390 20340 18510
rect 20220 18090 20340 18210
rect 23100 19290 23220 19410
rect 22860 18990 22980 19110
rect 23580 18990 23700 19110
rect 24810 19200 24930 19320
rect 25020 19170 25140 19290
rect 24540 18990 24660 19110
rect 25530 19170 25650 19290
rect 25740 19200 25860 19320
rect 25980 18990 26100 19110
rect 24990 18660 25110 18780
rect 24060 18390 24180 18510
rect 27420 19290 27540 19410
rect 24810 18360 24930 18480
rect 25740 18360 25860 18480
rect 26940 18390 27060 18510
rect 30540 18990 30660 19110
rect 31020 18390 31140 18510
rect 32460 18990 32580 19110
rect 33180 18990 33300 19110
rect 35580 18990 35700 19110
rect 35820 18990 35940 19110
rect 33420 18690 33540 18810
rect 32700 18390 32820 18510
rect 34860 18390 34980 18510
rect 37260 18990 37380 19110
rect 37980 18990 38100 19110
rect 36300 18390 36420 18510
rect 37500 18690 37620 18810
rect 37740 18090 37860 18210
rect 40620 19290 40740 19410
rect 40380 18990 40500 19110
rect 39420 18390 39540 18510
rect 39900 18390 40020 18510
rect 40860 18390 40980 18510
rect 45900 19590 46020 19710
rect 42060 18990 42180 19110
rect 43980 18990 44100 19110
rect 44460 18990 44580 19110
rect 42300 18690 42420 18810
rect 43740 18690 43860 18810
rect 44700 18690 44820 18810
rect 47340 18990 47460 19110
rect 48060 18990 48180 19110
rect 48060 18690 48180 18810
rect 49260 18690 49380 18810
rect 1214 17040 2086 17160
rect 53310 17040 54180 17160
rect 8010 15720 8130 15840
rect 8940 15720 9060 15840
rect 9690 15720 9810 15840
rect 10620 15720 10740 15840
rect 11310 15720 11430 15840
rect 12300 15720 12420 15840
rect 13470 15720 13590 15840
rect 14460 15720 14580 15840
rect 15210 15720 15330 15840
rect 16140 15720 16260 15840
rect 8190 15420 8310 15540
rect 9870 15420 9990 15540
rect 7740 15090 7860 15210
rect 6540 14790 6660 14910
rect 8010 14880 8130 15000
rect 8220 14910 8340 15030
rect 9180 15090 9300 15210
rect 9420 15090 9540 15210
rect 8730 14910 8850 15030
rect 8940 14880 9060 15000
rect 9690 14880 9810 15000
rect 9900 14910 10020 15030
rect 11700 15120 11820 15240
rect 10410 14910 10530 15030
rect 10620 14880 10740 15000
rect 11310 14880 11430 15000
rect 11580 14910 11700 15030
rect 15390 15420 15510 15540
rect 13020 15090 13140 15210
rect 13860 15120 13980 15240
rect 12090 14910 12210 15030
rect 12300 14880 12420 15000
rect 13470 14880 13590 15000
rect 13740 14910 13860 15030
rect 14700 15090 14820 15210
rect 14940 15090 15060 15210
rect 14250 14910 14370 15030
rect 14460 14880 14580 15000
rect 15210 14880 15330 15000
rect 15420 14910 15540 15030
rect 16860 15090 16980 15210
rect 15930 14910 16050 15030
rect 16140 14880 16260 15000
rect 17820 15690 17940 15810
rect 18540 15390 18660 15510
rect 19260 15090 19380 15210
rect 20460 15690 20580 15810
rect 19980 15390 20100 15510
rect 21660 15690 21780 15810
rect 24060 15690 24180 15810
rect 20700 15090 20820 15210
rect 21900 15090 22020 15210
rect 19500 14790 19620 14910
rect 25980 15720 26100 15840
rect 26910 15720 27030 15840
rect 26730 15420 26850 15540
rect 28380 15690 28500 15810
rect 25260 15090 25380 15210
rect 25500 15090 25620 15210
rect 25980 14880 26100 15000
rect 26190 14910 26310 15030
rect 21900 14490 22020 14610
rect 27900 15090 28020 15210
rect 26700 14910 26820 15030
rect 26910 14880 27030 15000
rect 28620 15390 28740 15510
rect 30540 15720 30660 15840
rect 31470 15720 31590 15840
rect 28380 15090 28500 15210
rect 29100 15090 29220 15210
rect 31290 15420 31410 15540
rect 30300 15090 30420 15210
rect 30540 14880 30660 15000
rect 30750 14910 30870 15030
rect 31740 15090 31860 15210
rect 31260 14910 31380 15030
rect 31470 14880 31590 15000
rect 32940 15090 33060 15210
rect 33180 15090 33300 15210
rect 33660 15690 33780 15810
rect 33660 15090 33780 15210
rect 34620 15090 34740 15210
rect 34380 14790 34500 14910
rect 35580 15690 35700 15810
rect 37740 15690 37860 15810
rect 37740 15090 37860 15210
rect 35820 14790 35940 14910
rect 38220 15690 38340 15810
rect 38940 15720 39060 15840
rect 39870 15720 39990 15840
rect 41850 15720 41970 15840
rect 42780 15720 42900 15840
rect 38700 15390 38820 15510
rect 39690 15420 39810 15540
rect 42030 15420 42150 15540
rect 38460 15090 38580 15210
rect 38940 14880 39060 15000
rect 39150 14910 39270 15030
rect 41340 15090 41460 15210
rect 41580 15090 41700 15210
rect 44700 15390 44820 15510
rect 39660 14910 39780 15030
rect 39870 14880 39990 15000
rect 41850 14880 41970 15000
rect 42060 14910 42180 15030
rect 43500 15090 43620 15210
rect 44460 15090 44580 15210
rect 45180 15090 45300 15210
rect 42570 14910 42690 15030
rect 42780 14880 42900 15000
rect 46860 15690 46980 15810
rect 49980 15690 50100 15810
rect 48060 15090 48180 15210
rect 48780 15090 48900 15210
rect 3194 14040 4066 14160
rect 51330 14040 52200 14160
rect 5580 13290 5700 13410
rect 11580 13590 11700 13710
rect 6540 12390 6660 12510
rect 7740 12990 7860 13110
rect 8460 12990 8580 13110
rect 9900 12990 10020 13110
rect 9180 12690 9300 12810
rect 9660 12690 9780 12810
rect 15900 12990 16020 13110
rect 11580 12390 11700 12510
rect 12540 12690 12660 12810
rect 17850 13200 17970 13320
rect 18060 13170 18180 13290
rect 17340 12990 17460 13110
rect 18570 13170 18690 13290
rect 18780 13200 18900 13320
rect 19500 13200 19620 13320
rect 16380 12390 16500 12510
rect 19710 13170 19830 13290
rect 17100 12690 17220 12810
rect 20220 13170 20340 13290
rect 20490 13200 20610 13320
rect 22110 13200 22230 13320
rect 22380 13170 22500 13290
rect 20100 12960 20220 13080
rect 18030 12660 18150 12780
rect 22500 12960 22620 13080
rect 22890 13170 23010 13290
rect 23100 13200 23220 13320
rect 25020 12990 25140 13110
rect 25500 12990 25620 13110
rect 28140 12990 28260 13110
rect 29100 12990 29220 13110
rect 29340 12690 29460 12810
rect 17850 12360 17970 12480
rect 18780 12360 18900 12480
rect 19500 12360 19620 12480
rect 20490 12360 20610 12480
rect 22110 12360 22230 12480
rect 23100 12360 23220 12480
rect 27900 12390 28020 12510
rect 30060 12390 30180 12510
rect 33210 13200 33330 13320
rect 33420 13170 33540 13290
rect 33930 13170 34050 13290
rect 34140 13200 34260 13320
rect 35580 12990 35700 13110
rect 33390 12660 33510 12780
rect 36540 12990 36660 13110
rect 37020 12990 37140 13110
rect 33210 12360 33330 12480
rect 34140 12360 34260 12480
rect 37980 12990 38100 13110
rect 38460 12990 38580 13110
rect 38700 12990 38820 13110
rect 39900 12990 40020 13110
rect 41100 12990 41220 13110
rect 41580 12990 41700 13110
rect 37980 12390 38100 12510
rect 39420 12390 39540 12510
rect 43260 12990 43380 13110
rect 43980 12990 44100 13110
rect 45180 12990 45300 13110
rect 43020 12090 43140 12210
rect 44700 12690 44820 12810
rect 43740 12390 43860 12510
rect 46620 12990 46740 13110
rect 47580 12990 47700 13110
rect 47820 12690 47940 12810
rect 49740 12990 49860 13110
rect 49020 12390 49140 12510
rect 49980 12690 50100 12810
rect 1214 11040 2086 11160
rect 53310 11040 54180 11160
rect 6300 9390 6420 9510
rect 5340 9090 5460 9210
rect 6780 9090 6900 9210
rect 7260 9690 7380 9810
rect 8010 9720 8130 9840
rect 8940 9720 9060 9840
rect 9420 10590 9540 10710
rect 8190 9420 8310 9540
rect 8010 8880 8130 9000
rect 8220 8910 8340 9030
rect 9420 9090 9540 9210
rect 8730 8910 8850 9030
rect 8940 8880 9060 9000
rect 10140 9690 10260 9810
rect 11100 9690 11220 9810
rect 10380 9090 10500 9210
rect 14010 9720 14130 9840
rect 14940 9720 15060 9840
rect 14190 9420 14310 9540
rect 12540 9090 12660 9210
rect 12780 9090 12900 9210
rect 14010 8880 14130 9000
rect 14220 8910 14340 9030
rect 15180 9090 15300 9210
rect 14730 8910 14850 9030
rect 14940 8880 15060 9000
rect 17100 9690 17220 9810
rect 17550 9720 17670 9840
rect 18540 9720 18660 9840
rect 19500 9720 19620 9840
rect 20430 9720 20550 9840
rect 20940 9690 21060 9810
rect 20250 9420 20370 9540
rect 17940 9120 18060 9240
rect 17550 8880 17670 9000
rect 17820 8910 17940 9030
rect 18330 8910 18450 9030
rect 18540 8880 18660 9000
rect 19500 8880 19620 9000
rect 19710 8910 19830 9030
rect 20700 9090 20820 9210
rect 21180 9090 21300 9210
rect 20220 8910 20340 9030
rect 20430 8880 20550 9000
rect 22140 9720 22260 9840
rect 23070 9720 23190 9840
rect 22890 9420 23010 9540
rect 21900 9090 22020 9210
rect 21420 8790 21540 8910
rect 22140 8880 22260 9000
rect 22350 8910 22470 9030
rect 23340 9090 23460 9210
rect 23820 9090 23940 9210
rect 22860 8910 22980 9030
rect 23070 8880 23190 9000
rect 24540 9690 24660 9810
rect 25260 9690 25380 9810
rect 25770 9720 25890 9840
rect 26700 9720 26820 9840
rect 25950 9420 26070 9540
rect 24300 9090 24420 9210
rect 25020 9090 25140 9210
rect 25770 8880 25890 9000
rect 25980 8910 26100 9030
rect 26940 9090 27060 9210
rect 27420 9090 27540 9210
rect 26490 8910 26610 9030
rect 26700 8880 26820 9000
rect 28380 9690 28500 9810
rect 28860 9690 28980 9810
rect 29580 8790 29700 8910
rect 32460 9690 32580 9810
rect 33420 9720 33540 9840
rect 34410 9720 34530 9840
rect 35580 9990 35700 10110
rect 31740 9090 31860 9210
rect 32220 9090 32340 9210
rect 33180 9090 33300 9210
rect 33420 8880 33540 9000
rect 33630 8910 33750 9030
rect 34020 9120 34140 9240
rect 35340 9090 35460 9210
rect 34140 8910 34260 9030
rect 34410 8880 34530 9000
rect 36300 9090 36420 9210
rect 37260 9690 37380 9810
rect 38460 9090 38580 9210
rect 38940 9090 39060 9210
rect 39900 9090 40020 9210
rect 40860 9690 40980 9810
rect 41100 9090 41220 9210
rect 42810 9720 42930 9840
rect 43740 9720 43860 9840
rect 45450 9720 45570 9840
rect 46380 9720 46500 9840
rect 42990 9420 43110 9540
rect 43980 9390 44100 9510
rect 44460 9390 44580 9510
rect 45630 9420 45750 9540
rect 47580 9690 47700 9810
rect 47580 9390 47700 9510
rect 42540 9090 42660 9210
rect 42810 8880 42930 9000
rect 43020 8910 43140 9030
rect 45180 9090 45300 9210
rect 43530 8910 43650 9030
rect 43740 8880 43860 9000
rect 45450 8880 45570 9000
rect 45660 8910 45780 9030
rect 46860 9090 46980 9210
rect 46170 8910 46290 9030
rect 46380 8880 46500 9000
rect 48300 9090 48420 9210
rect 3194 8040 4066 8160
rect 51330 8040 52200 8160
rect 5820 7200 5940 7320
rect 6030 7170 6150 7290
rect 7260 7590 7380 7710
rect 6540 7170 6660 7290
rect 6750 7200 6870 7320
rect 7740 6990 7860 7110
rect 6570 6660 6690 6780
rect 5820 6360 5940 6480
rect 6750 6360 6870 6480
rect 8460 6990 8580 7110
rect 9900 6990 10020 7110
rect 8220 6390 8340 6510
rect 9420 6690 9540 6810
rect 12300 6690 12420 6810
rect 13020 6990 13140 7110
rect 15420 7290 15540 7410
rect 15900 7290 16020 7410
rect 16860 7290 16980 7410
rect 20940 7290 21060 7410
rect 12780 6690 12900 6810
rect 18540 6990 18660 7110
rect 20700 6990 20820 7110
rect 18540 6690 18660 6810
rect 21180 6990 21300 7110
rect 23340 6990 23460 7110
rect 21420 6390 21540 6510
rect 24300 7290 24420 7410
rect 25950 7200 26070 7320
rect 26220 7170 26340 7290
rect 26340 6960 26460 7080
rect 26730 7170 26850 7290
rect 26940 7200 27060 7320
rect 28140 7290 28260 7410
rect 27660 6990 27780 7110
rect 27900 6690 28020 6810
rect 25260 6390 25380 6510
rect 25950 6360 26070 6480
rect 26940 6360 27060 6480
rect 28380 6990 28500 7110
rect 30330 7200 30450 7320
rect 30540 7170 30660 7290
rect 36780 7590 36900 7710
rect 31050 7170 31170 7290
rect 31260 7200 31380 7320
rect 32460 6990 32580 7110
rect 30510 6660 30630 6780
rect 29580 6390 29700 6510
rect 30330 6360 30450 6480
rect 31260 6360 31380 6480
rect 33660 6390 33780 6510
rect 35100 6990 35220 7110
rect 35340 6990 35460 7110
rect 38700 6990 38820 7110
rect 36540 6390 36660 6510
rect 39420 6990 39540 7110
rect 39660 6990 39780 7110
rect 42540 7290 42660 7410
rect 42060 6990 42180 7110
rect 42540 6990 42660 7110
rect 44220 6990 44340 7110
rect 40860 6390 40980 6510
rect 43980 6690 44100 6810
rect 44460 6690 44580 6810
rect 48060 6990 48180 7110
rect 47340 6390 47460 6510
rect 47820 6690 47940 6810
rect 1214 5040 2086 5160
rect 53310 5040 54180 5160
rect 3194 3104 4066 3976
rect 51330 3104 52200 3976
rect 17100 2790 17220 2910
rect 35580 2790 35700 2910
rect 17340 2490 17460 2610
rect 28620 2490 28740 2610
rect 18540 2190 18660 2310
rect 21180 2190 21300 2310
rect 1214 1124 2086 1996
rect 53310 1124 54180 1996
<< metal2 >>
rect 1155 48076 2145 48135
rect 1155 47204 1214 48076
rect 2086 47204 2145 48076
rect 1155 41160 2145 47204
rect 1155 41040 1214 41160
rect 2086 41040 2145 41160
rect 1155 35160 2145 41040
rect 3135 46096 4125 46155
rect 3135 45224 3194 46096
rect 4066 45224 4125 46096
rect 3135 44160 4125 45224
rect 3135 44040 3194 44160
rect 4066 44040 4125 44160
rect 1155 35040 1214 35160
rect 2086 35040 2145 35160
rect 1155 29160 2145 35040
rect 1155 29040 1214 29160
rect 2086 29040 2145 29160
rect 795 0 885 26190
rect 1155 23160 2145 29040
rect 1155 23040 1214 23160
rect 2086 23040 2145 23160
rect 1155 17160 2145 23040
rect 1155 17040 1214 17160
rect 2086 17040 2145 17160
rect 1155 11160 2145 17040
rect 2475 16110 2565 38790
rect 3135 38160 4125 44040
rect 9435 44010 9525 49200
rect 14475 49110 14565 49200
rect 14460 48990 14580 49110
rect 9330 43200 9420 43290
rect 5355 38160 5445 42990
rect 7275 42510 7365 42990
rect 8715 42810 8805 42990
rect 8955 42510 9045 42990
rect 9210 42480 9300 43200
rect 9540 43200 9930 43290
rect 10170 43080 10260 43200
rect 12795 43110 12885 43290
rect 9420 42990 10260 43080
rect 9420 42780 9510 42990
rect 7275 40710 7365 42390
rect 8475 40710 8565 42390
rect 10170 42480 10260 42990
rect 8460 40590 8580 40710
rect 9675 39510 9765 42390
rect 10395 41295 10485 42990
rect 10155 41205 10485 41295
rect 10155 39810 10245 41205
rect 10635 40995 10725 42990
rect 10875 42810 10965 42990
rect 10395 40905 10725 40995
rect 3135 38040 3194 38160
rect 4066 38040 4125 38160
rect 2820 37605 3045 37695
rect 2715 13410 2805 37290
rect 1155 11040 1214 11160
rect 2086 11040 2145 11160
rect 1155 5160 2145 11040
rect 2955 6495 3045 37605
rect 2820 6405 3045 6495
rect 3135 32160 4125 38040
rect 5595 36795 5685 39390
rect 9675 39210 9765 39390
rect 7035 37710 7125 38790
rect 7515 37710 7605 39090
rect 3135 32040 3194 32160
rect 4066 32040 4125 32160
rect 3135 26160 4125 32040
rect 5355 36705 5685 36795
rect 5355 31110 5445 36705
rect 5820 35490 5940 35610
rect 5835 33810 5925 35490
rect 7035 33510 7125 36390
rect 7275 33810 7365 36990
rect 6555 32760 6645 33090
rect 7035 31710 7125 33390
rect 7275 33210 7365 33690
rect 7515 33210 7605 37290
rect 8475 36195 8565 36990
rect 10155 36210 10245 39690
rect 10395 38910 10485 40905
rect 11355 39510 11445 39990
rect 11595 39210 11685 42690
rect 12795 40110 12885 42990
rect 13035 42810 13125 43290
rect 11790 39000 11880 39720
rect 12810 39210 12900 39720
rect 12300 39120 12900 39210
rect 12180 38910 12570 39000
rect 12810 39000 12900 39120
rect 10860 38490 10980 38610
rect 10875 37410 10965 38490
rect 12075 37710 12165 38910
rect 12300 38490 12420 38610
rect 12315 37710 12405 38490
rect 13515 37710 13605 39090
rect 12060 37590 12180 37710
rect 11355 36510 11445 36690
rect 12075 36510 12165 37290
rect 13035 36510 13125 36990
rect 8235 36105 8565 36195
rect 5580 31080 5670 31200
rect 5910 31200 6300 31290
rect 5580 30990 6180 31080
rect 5355 30510 5445 30990
rect 5580 30480 5670 30990
rect 6600 30480 6690 31200
rect 3135 26040 3194 26160
rect 4066 26040 4125 26160
rect 3135 20160 4125 26040
rect 6075 25710 6165 27240
rect 7035 27210 7125 30990
rect 7290 27000 7380 27720
rect 7755 27510 7845 33690
rect 8235 33510 8325 36105
rect 11835 34710 11925 36390
rect 11820 34590 11940 34710
rect 8235 31410 8325 33390
rect 8715 31710 8805 33090
rect 9150 33000 9240 33720
rect 10170 33210 10260 33720
rect 9660 33120 10260 33210
rect 9540 32910 9930 33000
rect 10170 33000 10260 33120
rect 8700 31590 8820 31710
rect 8235 28995 8325 30690
rect 8475 30510 8565 30990
rect 9195 30510 9285 30990
rect 8235 28905 8565 28995
rect 7500 27210 7590 27420
rect 8250 27210 8340 27720
rect 8475 27210 8565 28905
rect 8955 28710 9045 30390
rect 9435 30210 9525 32910
rect 9660 32490 9780 32610
rect 9675 31110 9765 32490
rect 10875 32310 10965 33090
rect 11310 33000 11400 33720
rect 12330 33210 12420 33720
rect 11820 33120 12420 33210
rect 11700 32910 12090 33000
rect 12330 33000 12420 33120
rect 11835 31710 11925 32190
rect 11820 31590 11940 31710
rect 11490 31200 11580 31290
rect 10155 30810 10245 30990
rect 8940 28590 9060 28710
rect 9195 27810 9285 29490
rect 9195 27210 9285 27390
rect 9660 27210 9750 27720
rect 7500 27120 8340 27210
rect 7410 26910 7500 27000
rect 7620 26910 8010 27000
rect 8250 27000 8340 27120
rect 9660 27120 10260 27210
rect 8715 26910 8805 27090
rect 9660 27000 9750 27120
rect 9990 26910 10380 27000
rect 10680 27000 10770 27720
rect 11115 27210 11205 30990
rect 11370 30480 11460 31200
rect 11700 31200 12090 31290
rect 12330 31080 12420 31200
rect 12795 31110 12885 33990
rect 11580 30990 12420 31080
rect 11580 30780 11670 30990
rect 12330 30480 12420 30990
rect 11355 27510 11445 27690
rect 11835 27210 11925 30390
rect 12075 29910 12165 30090
rect 12075 27210 12165 29790
rect 12555 27210 12645 27990
rect 12795 27810 12885 30990
rect 13035 30510 13125 36390
rect 13755 34710 13845 36690
rect 13740 34590 13860 34710
rect 13995 34110 14085 39690
rect 14235 39210 14325 42990
rect 14475 40710 14565 48990
rect 14460 40590 14580 40710
rect 13995 31110 14085 32790
rect 13755 28710 13845 30690
rect 13740 28590 13860 28710
rect 14475 28110 14565 39990
rect 15195 39210 15285 46590
rect 18075 45195 18165 46890
rect 17835 45105 18165 45195
rect 17115 43110 17205 43290
rect 15915 42510 16005 42690
rect 15675 39810 15765 41190
rect 17595 39810 17685 42990
rect 14955 32910 15045 36390
rect 15195 34410 15285 39090
rect 15435 37110 15525 38790
rect 16155 38610 16245 39090
rect 17100 38490 17220 38610
rect 15675 33810 15765 36690
rect 15675 32910 15765 33690
rect 15915 33210 16005 36990
rect 16155 36510 16245 38490
rect 17115 37410 17205 38490
rect 17355 38295 17445 39690
rect 17595 38610 17685 38790
rect 17580 38490 17700 38610
rect 17355 38205 17685 38295
rect 17595 37110 17685 38205
rect 16395 33210 16485 36990
rect 14910 30480 15000 31200
rect 15300 31200 15690 31290
rect 15930 31080 16020 31200
rect 15420 30990 16020 31080
rect 15930 30480 16020 30990
rect 15420 29490 15540 29610
rect 15435 27510 15525 29490
rect 16395 27810 16485 32490
rect 16635 30795 16725 33090
rect 17115 32610 17205 36390
rect 17355 33810 17445 36990
rect 17595 33510 17685 36990
rect 17835 36510 17925 45105
rect 18555 43710 18645 49200
rect 18075 42510 18165 42690
rect 18795 39510 18885 42390
rect 19035 38910 19125 43290
rect 19500 43080 19590 43200
rect 19830 43200 20220 43290
rect 19500 42990 20100 43080
rect 19275 42510 19365 42990
rect 19500 42480 19590 42990
rect 20520 42480 20610 43200
rect 19755 39210 19845 42390
rect 20955 39810 21045 43290
rect 22395 40695 22485 43890
rect 27675 43710 27765 49200
rect 31515 43410 31605 43590
rect 23010 43200 23100 43290
rect 22635 41010 22725 42990
rect 22890 42480 22980 43200
rect 23220 43200 23610 43290
rect 23850 43080 23940 43200
rect 23100 42990 23940 43080
rect 23100 42780 23190 42990
rect 23850 42480 23940 42990
rect 25755 42210 25845 42990
rect 27195 42795 27285 42990
rect 26955 42705 27285 42795
rect 22620 40695 22740 40710
rect 22395 40605 22740 40695
rect 22620 40590 22740 40605
rect 20955 39210 21045 39690
rect 21435 39210 21525 39390
rect 21060 39105 21285 39195
rect 18555 36510 18645 36990
rect 18300 35490 18420 35610
rect 18315 33810 18405 35490
rect 17340 32490 17460 32610
rect 17355 31710 17445 32490
rect 16875 31110 16965 31590
rect 16635 30705 16965 30795
rect 16875 28710 16965 30705
rect 17115 30210 17205 30990
rect 17310 30480 17400 31200
rect 17700 31200 18090 31290
rect 18330 31080 18420 31200
rect 17820 30990 18420 31080
rect 18330 30480 18420 30990
rect 16860 28590 16980 28710
rect 10140 26490 10260 26610
rect 7755 25710 7845 26490
rect 10155 26010 10245 26490
rect 6060 25590 6180 25710
rect 7740 25590 7860 25710
rect 9435 25410 9525 25890
rect 5730 25200 5820 25290
rect 5610 24480 5700 25200
rect 5940 25200 6330 25290
rect 6570 25080 6660 25200
rect 8475 25110 8565 25290
rect 9435 25110 9525 25290
rect 9810 25200 9900 25290
rect 5820 24990 6660 25080
rect 5820 24780 5910 24990
rect 6570 24480 6660 24990
rect 6795 24810 6885 24990
rect 3135 20040 3194 20160
rect 4066 20040 4125 20160
rect 3135 14160 4125 20040
rect 5355 19710 5445 21090
rect 5610 21000 5700 21720
rect 5820 21210 5910 21420
rect 6570 21210 6660 21720
rect 7035 21510 7125 24990
rect 9195 24510 9285 24990
rect 9690 24480 9780 25200
rect 10020 25200 10410 25290
rect 10650 25080 10740 25200
rect 9900 24990 10740 25080
rect 9900 24780 9990 24990
rect 10650 24480 10740 24990
rect 9675 21510 9765 21690
rect 10155 21210 10245 21690
rect 10395 21210 10485 21390
rect 5820 21120 6660 21210
rect 5730 20910 5820 21000
rect 5940 20910 6330 21000
rect 6570 21000 6660 21120
rect 6795 20910 6885 21090
rect 8955 20610 9045 21090
rect 8955 19110 9045 20490
rect 9675 19710 9765 20790
rect 9660 19590 9780 19710
rect 10155 19695 10245 21090
rect 11595 20610 11685 21390
rect 10155 19605 10485 19695
rect 9180 19080 9270 19200
rect 9510 19200 9900 19290
rect 10020 19200 10110 19290
rect 9180 18990 10020 19080
rect 3135 14040 3194 14160
rect 4066 14040 4125 14160
rect 3135 8160 4125 14040
rect 5595 13410 5685 18390
rect 6075 15210 6165 18690
rect 6795 15810 6885 18990
rect 9180 18480 9270 18990
rect 9930 18780 10020 18990
rect 10140 18480 10230 19200
rect 10395 19110 10485 19605
rect 9435 15810 9525 16290
rect 6555 12510 6645 14790
rect 5355 9210 5445 11040
rect 6315 9510 6405 9990
rect 6795 9210 6885 9390
rect 3135 8040 3194 8160
rect 4066 8040 4125 8160
rect 1155 5040 1214 5160
rect 2086 5040 2145 5160
rect 1155 1996 2145 5040
rect 3135 3976 4125 8040
rect 5820 7080 5910 7200
rect 6150 7200 6540 7290
rect 6660 7200 6750 7290
rect 5820 6990 6660 7080
rect 5820 6480 5910 6990
rect 6570 6780 6660 6990
rect 6780 6480 6870 7200
rect 7035 6210 7125 13590
rect 7755 13110 7845 15090
rect 8010 15000 8100 15720
rect 8220 15210 8310 15420
rect 8970 15210 9060 15720
rect 9195 15210 9285 15390
rect 9435 15210 9525 15690
rect 8220 15120 9060 15210
rect 8130 14910 8220 15000
rect 8340 14910 8730 15000
rect 8970 15000 9060 15120
rect 9690 15000 9780 15720
rect 9900 15210 9990 15420
rect 10650 15210 10740 15720
rect 10875 15210 10965 17490
rect 9900 15120 10740 15210
rect 9810 14910 9900 15000
rect 10020 14910 10410 15000
rect 10650 15000 10740 15120
rect 8475 10110 8565 12990
rect 9675 12810 9765 14490
rect 11115 14310 11205 18990
rect 11595 18510 11685 20490
rect 12075 19290 12165 23490
rect 12315 19710 12405 21090
rect 12300 19590 12420 19710
rect 13275 19695 13365 27390
rect 16635 27210 16725 27690
rect 15195 26610 15285 27090
rect 15435 26310 15525 27090
rect 17595 26010 17685 30090
rect 18795 27810 18885 34290
rect 19035 33210 19125 38790
rect 21195 37410 21285 39105
rect 19515 36810 19605 36990
rect 19995 33210 20085 36390
rect 21435 36210 21525 36390
rect 21195 32910 21285 33690
rect 21675 32310 21765 39090
rect 21915 38910 22005 39090
rect 22170 39000 22260 39720
rect 22380 39210 22470 39420
rect 23130 39210 23220 39720
rect 24075 39510 24165 40890
rect 25755 39810 25845 42090
rect 26235 40710 26325 42690
rect 26955 40710 27045 42705
rect 27915 42510 28005 42990
rect 28155 42810 28245 42990
rect 29595 42510 29685 42990
rect 31275 42810 31365 42990
rect 27195 42210 27285 42390
rect 26940 40590 27060 40710
rect 24075 39210 24165 39390
rect 24315 39210 24405 39390
rect 22380 39120 23220 39210
rect 22290 38910 22380 39000
rect 22500 38910 22890 39000
rect 23130 39000 23220 39120
rect 24795 38910 24885 39090
rect 25755 38910 25845 39690
rect 26235 39510 26325 40590
rect 22395 37110 22485 37290
rect 23835 37110 23925 37290
rect 22875 35910 22965 36390
rect 22620 35490 22740 35610
rect 22635 33210 22725 35490
rect 22875 33510 22965 35790
rect 19275 31110 19365 31290
rect 19650 31200 19740 31290
rect 19035 30810 19125 30990
rect 19530 30480 19620 31200
rect 19860 31200 20250 31290
rect 20490 31080 20580 31200
rect 21195 31110 21285 31290
rect 22875 31110 22965 31290
rect 19740 30990 20580 31080
rect 19740 30780 19830 30990
rect 20490 30480 20580 30990
rect 21675 30510 21765 30990
rect 17835 27210 17925 27690
rect 19275 27510 19365 27690
rect 19755 27510 19845 29490
rect 13995 23610 14085 24390
rect 14235 22710 14325 24990
rect 15435 24810 15525 24990
rect 15675 24810 15765 24990
rect 14235 21210 14325 22590
rect 14490 21000 14580 21720
rect 14700 21210 14790 21420
rect 15450 21210 15540 21720
rect 15675 21210 15765 24690
rect 14700 21120 15540 21210
rect 14610 20910 14700 21000
rect 14820 20910 15210 21000
rect 15450 21000 15540 21120
rect 14940 20490 15060 20610
rect 13035 19605 13365 19695
rect 11790 18480 11880 19200
rect 12180 19200 12570 19290
rect 12810 19080 12900 19200
rect 12300 18990 12900 19080
rect 12810 18480 12900 18990
rect 13035 18795 13125 19605
rect 14955 19410 15045 20490
rect 15675 20310 15765 21090
rect 16875 19410 16965 20490
rect 13275 19110 13365 19290
rect 13890 19200 13980 19290
rect 13515 18810 13605 18990
rect 13035 18705 13365 18795
rect 11310 15000 11400 15720
rect 12330 15210 12420 15720
rect 11820 15120 12420 15210
rect 11700 14910 12090 15000
rect 12330 15000 12420 15120
rect 12555 14910 12645 15990
rect 13035 15210 13125 15690
rect 11595 13710 11685 14190
rect 9915 13110 10005 13290
rect 12795 13110 12885 14190
rect 9195 11295 9285 12690
rect 9195 11205 9525 11295
rect 9435 10710 9525 11205
rect 7275 9810 7365 9990
rect 7275 7710 7365 9690
rect 8010 9000 8100 9720
rect 8220 9210 8310 9420
rect 8970 9210 9060 9720
rect 9435 9210 9525 9390
rect 9675 9210 9765 12690
rect 9915 9510 10005 12990
rect 12555 12510 12645 12690
rect 11100 11490 11220 11610
rect 11115 9810 11205 11490
rect 11595 10710 11685 12390
rect 11580 10590 11700 10710
rect 10155 9210 10245 9690
rect 10395 9210 10485 9390
rect 12555 9210 12645 9690
rect 12795 9210 12885 12990
rect 8220 9120 9060 9210
rect 8130 8910 8220 9000
rect 8340 8910 8730 9000
rect 8970 9000 9060 9120
rect 7755 6210 7845 6990
rect 8235 6510 8325 7290
rect 6300 5490 6420 5610
rect 3135 3104 3194 3976
rect 4066 3104 4125 3976
rect 3135 3045 4125 3104
rect 1155 1124 1214 1996
rect 2086 1124 2145 1996
rect 1155 1065 2145 1124
rect 6315 840 6405 5490
rect 6555 0 6645 6090
rect 8475 5760 8565 6990
rect 9915 6810 10005 6990
rect 12795 6810 12885 6990
rect 9435 6510 9525 6690
rect 12315 6510 12405 6690
rect 13035 6210 13125 6990
rect 13275 6510 13365 18705
rect 13770 18480 13860 19200
rect 14100 19200 14490 19290
rect 14730 19080 14820 19200
rect 13980 18990 14820 19080
rect 13980 18780 14070 18990
rect 14730 18480 14820 18990
rect 15675 18810 15765 18990
rect 14220 17490 14340 17610
rect 14235 15810 14325 17490
rect 16395 16110 16485 18390
rect 13470 15000 13560 15720
rect 14490 15210 14580 15720
rect 14715 15210 14805 15390
rect 14955 15210 15045 15690
rect 13980 15120 14580 15210
rect 13860 14910 14250 15000
rect 14490 15000 14580 15120
rect 15210 15000 15300 15720
rect 15420 15210 15510 15420
rect 16170 15210 16260 15720
rect 16875 15210 16965 15690
rect 15420 15120 16260 15210
rect 15330 14910 15420 15000
rect 15540 14910 15930 15000
rect 16170 15000 16260 15120
rect 17115 14610 17205 25890
rect 18075 23010 18165 27090
rect 18075 21210 18165 22290
rect 18315 21210 18405 26790
rect 18795 26610 18885 26790
rect 19755 24510 19845 27390
rect 20955 27210 21045 30090
rect 21195 28710 21285 30390
rect 22155 29910 22245 30990
rect 22635 30810 22725 30990
rect 21420 29490 21540 29610
rect 21180 28590 21300 28710
rect 21435 27810 21525 29490
rect 22875 28110 22965 30990
rect 23115 28110 23205 36090
rect 24060 35490 24180 35610
rect 24075 33510 24165 35490
rect 24315 33495 24405 37290
rect 24795 34410 24885 38790
rect 25035 36510 25125 36990
rect 25515 36810 25605 36990
rect 27195 36810 27285 39090
rect 25515 33810 25605 36690
rect 24315 33405 24645 33495
rect 23355 27795 23445 33390
rect 23595 31710 23685 33390
rect 24315 31410 24405 33090
rect 24075 30210 24165 30990
rect 23595 27810 23685 27990
rect 23115 27705 23445 27795
rect 21675 27210 21765 27690
rect 23115 27210 23205 27705
rect 24555 27510 24645 33405
rect 25275 33210 25365 33690
rect 25275 30510 25365 32790
rect 25515 31410 25605 33690
rect 25755 31710 25845 33090
rect 26250 33000 26340 33720
rect 26460 33210 26550 33420
rect 27210 33210 27300 33720
rect 27435 33210 27525 36990
rect 28875 36510 28965 41190
rect 29595 39810 29685 42390
rect 31275 42210 31365 42690
rect 31275 39210 31365 42090
rect 32235 40710 32325 42390
rect 32220 40590 32340 40710
rect 32475 39210 32565 42690
rect 32955 41895 33045 46590
rect 36555 43710 36645 49200
rect 45675 43710 45765 49200
rect 53250 48076 54240 48135
rect 53250 47204 53310 48076
rect 54180 47204 54240 48076
rect 51270 46096 52260 46155
rect 51270 45224 51330 46096
rect 52200 45224 52260 46096
rect 51270 44160 52260 45224
rect 51270 44040 51330 44160
rect 52200 44040 52260 44160
rect 34635 43110 34725 43290
rect 36210 43200 36300 43290
rect 33675 42810 33765 42990
rect 33195 42210 33285 42390
rect 32955 41805 33285 41895
rect 30795 37710 30885 38490
rect 31275 37710 31365 39090
rect 30780 37590 30900 37710
rect 32955 37410 33045 37590
rect 30075 37110 30165 37290
rect 28875 36210 28965 36390
rect 28395 35310 28485 36090
rect 26460 33120 27300 33210
rect 26370 32910 26460 33000
rect 26580 32910 26970 33000
rect 27210 33000 27300 33120
rect 29115 32910 29205 36990
rect 29595 35910 29685 36390
rect 30315 34710 30405 36690
rect 30300 34590 30420 34710
rect 30555 32910 30645 33990
rect 31035 33810 31125 37290
rect 32715 37110 32805 37290
rect 31755 36510 31845 36990
rect 31035 33510 31125 33690
rect 31995 33510 32085 36390
rect 32715 34110 32805 36990
rect 31515 33210 31605 33390
rect 31755 33210 31845 33390
rect 32955 33210 33045 36990
rect 33195 36510 33285 41805
rect 33690 39000 33780 39720
rect 33900 39210 33990 39420
rect 34650 39210 34740 39720
rect 35115 39210 35205 42990
rect 35355 39510 35445 42690
rect 33900 39120 34740 39210
rect 33810 38910 33900 39000
rect 34020 38910 34410 39000
rect 34650 39000 34740 39120
rect 33435 34710 33525 38790
rect 34875 37410 34965 39090
rect 34395 36510 34485 36990
rect 33420 34590 33540 34710
rect 25755 30810 25845 30990
rect 25995 30510 26085 30990
rect 25515 28110 25605 29490
rect 25515 27810 25605 27990
rect 21195 25110 21285 27090
rect 23355 25410 23445 27390
rect 25515 27210 25605 27390
rect 18555 21810 18645 22890
rect 17355 16710 17445 18390
rect 17340 16590 17460 16710
rect 16635 13710 16725 14490
rect 17595 14010 17685 21090
rect 17835 19710 17925 20790
rect 17820 19590 17940 19710
rect 17835 14910 17925 15690
rect 16620 13590 16740 13710
rect 15915 13110 16005 13290
rect 15195 10710 15285 12390
rect 16395 11295 16485 12390
rect 16395 11205 16725 11295
rect 16635 10710 16725 11205
rect 16620 10590 16740 10710
rect 14010 9000 14100 9720
rect 14220 9210 14310 9420
rect 14970 9210 15060 9720
rect 15195 9210 15285 10590
rect 14220 9120 15060 9210
rect 14130 8910 14220 9000
rect 14340 8910 14730 9000
rect 14970 9000 15060 9120
rect 16875 7410 16965 13890
rect 18075 13710 18165 21090
rect 18555 20910 18645 21690
rect 18795 21210 18885 24390
rect 19755 22410 19845 23490
rect 21195 23010 21285 24990
rect 19020 21210 19110 21720
rect 19770 21210 19860 21420
rect 19020 21120 19860 21210
rect 19020 21000 19110 21120
rect 19350 20910 19740 21000
rect 19980 21000 20070 21720
rect 20235 21210 20325 22890
rect 20700 21210 20790 21720
rect 21450 21210 21540 21420
rect 20700 21120 21540 21210
rect 19860 20910 19950 21000
rect 18315 19995 18405 20790
rect 18315 19905 18645 19995
rect 18555 19110 18645 19905
rect 19755 19410 19845 20190
rect 18315 17610 18405 18690
rect 19515 17910 19605 18990
rect 20235 18510 20325 20790
rect 20475 20610 20565 21090
rect 20700 21000 20790 21120
rect 21030 20910 21420 21000
rect 21660 21000 21750 21720
rect 21915 21210 22005 24990
rect 22155 21510 22245 21690
rect 22395 21210 22485 24990
rect 23595 24810 23685 27090
rect 24075 26610 24165 27090
rect 24075 25095 24165 26490
rect 25515 26010 25605 27090
rect 25755 26610 25845 30390
rect 23835 25005 24165 25095
rect 22635 21510 22725 21690
rect 21540 20910 21630 21000
rect 20955 18810 21045 18990
rect 18555 15510 18645 15690
rect 17970 13200 18060 13290
rect 17115 12810 17205 12990
rect 17115 9810 17205 12690
rect 15435 6510 15525 7290
rect 15915 7110 16005 7290
rect 17115 2910 17205 9690
rect 17355 9210 17445 12990
rect 17850 12480 17940 13200
rect 18180 13200 18570 13290
rect 18810 13080 18900 13200
rect 18060 12990 18900 13080
rect 18060 12780 18150 12990
rect 18810 12480 18900 12990
rect 17355 2610 17445 9090
rect 17550 9000 17640 9720
rect 18570 9210 18660 9720
rect 18060 9120 18660 9210
rect 17940 8910 18330 9000
rect 18570 9000 18660 9120
rect 17835 7710 17925 8910
rect 18795 8610 18885 9990
rect 19035 8910 19125 12690
rect 19275 10110 19365 15090
rect 19515 14310 19605 14790
rect 19995 13710 20085 15390
rect 20235 15210 20325 18090
rect 20475 15810 20565 15990
rect 19980 13590 20100 13710
rect 20235 13410 20325 13590
rect 19500 13080 19590 13200
rect 19830 13200 20220 13290
rect 19500 12990 20100 13080
rect 19500 12480 19590 12990
rect 20520 12480 20610 13200
rect 19980 11490 20100 11610
rect 19995 11010 20085 11490
rect 19500 9210 19590 9720
rect 20250 9210 20340 9420
rect 19500 9120 20340 9210
rect 19500 9000 19590 9120
rect 19830 8910 20220 9000
rect 20460 9000 20550 9720
rect 20715 9210 20805 15090
rect 21435 12510 21525 15690
rect 21675 12810 21765 15690
rect 21915 15210 22005 21090
rect 22635 19110 22725 21390
rect 23115 19410 23205 21390
rect 22875 18810 22965 18990
rect 23595 17010 23685 18990
rect 21915 14610 22005 14790
rect 22635 13710 22725 15390
rect 22620 13590 22740 13710
rect 22110 12480 22200 13200
rect 22500 13200 22890 13290
rect 23130 13080 23220 13200
rect 22620 12990 23220 13080
rect 23130 12480 23220 12990
rect 20955 9810 21045 10890
rect 22635 10710 22725 12390
rect 22620 10590 22740 10710
rect 20955 9210 21045 9690
rect 21915 9210 22005 9390
rect 22140 9210 22230 9720
rect 22890 9210 22980 9420
rect 21300 9105 21660 9195
rect 22140 9120 22980 9210
rect 20340 8910 20430 9000
rect 22140 9000 22230 9120
rect 22470 8910 22860 9000
rect 23100 9000 23190 9720
rect 23355 9210 23445 9690
rect 23835 9210 23925 25005
rect 24555 23910 24645 24690
rect 24075 18510 24165 19890
rect 24315 19110 24405 20790
rect 24555 20010 24645 23790
rect 25515 23610 25605 25890
rect 26235 25710 26325 32190
rect 31515 31710 31605 33090
rect 31500 31590 31620 31710
rect 33435 31410 33525 34290
rect 33675 33810 33765 36390
rect 34635 33795 34725 36990
rect 35115 36210 35205 36390
rect 35115 34110 35205 36090
rect 34635 33705 34965 33795
rect 26715 30510 26805 30990
rect 26715 28710 26805 30390
rect 26955 29310 27045 31290
rect 26700 28590 26820 28710
rect 27195 27810 27285 30690
rect 28395 29910 28485 30990
rect 28635 30510 28725 31290
rect 29835 31110 29925 31290
rect 31020 31080 31110 31200
rect 31350 31200 31740 31290
rect 31860 31200 31950 31290
rect 31020 30990 31860 31080
rect 27900 29490 28020 29610
rect 26220 25590 26340 25710
rect 25740 25080 25830 25200
rect 26070 25200 26460 25290
rect 26580 25200 26670 25290
rect 25740 24990 26580 25080
rect 25740 24480 25830 24990
rect 26490 24780 26580 24990
rect 26700 24480 26790 25200
rect 27195 24810 27285 27690
rect 25995 20010 26085 21690
rect 27435 21210 27525 24990
rect 26220 20490 26340 20610
rect 24555 19110 24645 19590
rect 26235 19410 26325 20490
rect 27435 19410 27525 21090
rect 24930 19200 25020 19290
rect 24075 16710 24165 18390
rect 24075 15510 24165 15690
rect 24315 11910 24405 16890
rect 24555 16110 24645 18990
rect 24810 18480 24900 19200
rect 25140 19200 25530 19290
rect 25770 19080 25860 19200
rect 25020 18990 25860 19080
rect 25020 18780 25110 18990
rect 25770 18480 25860 18990
rect 25995 16710 26085 18990
rect 27195 18495 27285 19290
rect 27060 18405 27285 18495
rect 24795 15795 24885 16590
rect 24555 15705 24885 15795
rect 24555 9810 24645 15705
rect 25275 15210 25365 15990
rect 25515 15210 25605 15390
rect 25980 15210 26070 15720
rect 26730 15210 26820 15420
rect 25980 15120 26820 15210
rect 25980 15000 26070 15120
rect 26310 14910 26700 15000
rect 26940 15000 27030 15720
rect 26820 14910 26910 15000
rect 26715 13110 26805 13290
rect 22980 8910 23070 9000
rect 23835 8910 23925 9090
rect 18555 7110 18645 7590
rect 20955 7410 21045 8790
rect 21195 7110 21285 8490
rect 18555 6210 18645 6690
rect 20715 6210 20805 6990
rect 18555 5310 18645 6090
rect 21195 2310 21285 6990
rect 21435 6510 21525 8790
rect 24315 7410 24405 9090
rect 24315 7110 24405 7290
rect 23355 5910 23445 6990
rect 12540 870 12660 900
rect 12540 90 12660 750
rect 12555 0 12645 90
rect 18555 0 18645 2190
rect 24555 0 24645 8790
rect 24795 870 24885 11790
rect 25035 9210 25125 12990
rect 25515 9810 25605 12990
rect 26235 10710 26325 12990
rect 26220 10590 26340 10710
rect 25275 6510 25365 9690
rect 25770 9000 25860 9720
rect 25980 9210 26070 9420
rect 26730 9210 26820 9720
rect 26955 9210 27045 12690
rect 27435 9210 27525 18090
rect 27675 16410 27765 29490
rect 27915 27810 28005 29490
rect 28635 27210 28725 30090
rect 29115 29910 29205 30390
rect 30075 30210 30165 30990
rect 31020 30480 31110 30990
rect 31770 30780 31860 30990
rect 31980 30480 32070 31200
rect 32235 31110 32325 31290
rect 29115 27210 29205 29790
rect 33195 28110 33285 30990
rect 33675 30510 33765 33690
rect 34635 32910 34725 33090
rect 33915 29610 34005 30990
rect 33675 28710 33765 29190
rect 33660 28590 33780 28710
rect 27915 24510 28005 24990
rect 29115 23610 29205 27090
rect 29355 25110 29445 27690
rect 30315 27510 30405 27690
rect 30795 26910 30885 27090
rect 29355 24510 29445 24690
rect 30795 24510 30885 26790
rect 32235 26295 32325 27390
rect 32475 26910 32565 27090
rect 32235 26205 32565 26295
rect 32475 25410 32565 26205
rect 32715 25410 32805 27090
rect 31755 25110 31845 25290
rect 28155 21210 28245 23490
rect 28395 19710 28485 21390
rect 28380 19590 28500 19710
rect 29355 18795 29445 24390
rect 29595 19110 29685 21390
rect 29835 21210 29925 21690
rect 30795 21210 30885 24090
rect 30555 19110 30645 20490
rect 31035 20310 31125 24390
rect 31755 24210 31845 24990
rect 32475 24810 32565 25290
rect 32955 24210 33045 27690
rect 33210 27000 33300 27720
rect 33420 27210 33510 27420
rect 34170 27210 34260 27720
rect 34635 27210 34725 32790
rect 34875 29910 34965 33705
rect 35115 33210 35205 33690
rect 35355 33210 35445 35790
rect 35115 31710 35205 33090
rect 35115 31110 35205 31290
rect 35595 30210 35685 39090
rect 35835 37710 35925 42990
rect 36090 42480 36180 43200
rect 36420 43200 36810 43290
rect 37050 43080 37140 43200
rect 36300 42990 37140 43080
rect 39660 43080 39750 43200
rect 39990 43200 40380 43290
rect 40500 43200 40590 43290
rect 45540 43305 45765 43395
rect 39660 42990 40500 43080
rect 36300 42780 36390 42990
rect 37050 42480 37140 42990
rect 37275 39810 37365 42990
rect 37755 41295 37845 42390
rect 37755 41205 38085 41295
rect 37995 40710 38085 41205
rect 37980 40590 38100 40710
rect 37275 37410 37365 39690
rect 38235 39210 38325 42690
rect 38235 38910 38325 39090
rect 35820 37080 35910 37200
rect 36150 37200 36540 37290
rect 36660 37200 36750 37290
rect 35820 36990 36660 37080
rect 35820 36480 35910 36990
rect 36570 36780 36660 36990
rect 36780 36480 36870 37200
rect 37035 37110 37125 37290
rect 36315 34710 36405 34890
rect 36300 34590 36420 34710
rect 35835 31410 35925 33090
rect 36315 30810 36405 33990
rect 37035 32610 37125 36990
rect 37275 34710 37365 37290
rect 38715 34110 38805 39390
rect 39435 39210 39525 42990
rect 39660 42480 39750 42990
rect 40410 42780 40500 42990
rect 40620 42480 40710 43200
rect 40875 43110 40965 43290
rect 40875 39510 40965 39690
rect 42315 39510 42405 42990
rect 41595 38910 41685 39390
rect 42555 39210 42645 43290
rect 45060 43005 45285 43095
rect 40470 37590 40500 37710
rect 39435 36810 39525 37590
rect 40395 37410 40485 37590
rect 40635 37110 40725 38490
rect 40875 36810 40965 38790
rect 39435 33810 39525 36390
rect 39435 33510 39525 33690
rect 40395 33510 40485 35490
rect 40875 33510 40965 36690
rect 35115 28710 35205 30090
rect 35100 28590 35220 28710
rect 33420 27120 34260 27210
rect 33330 26910 33420 27000
rect 33540 26910 33930 27000
rect 34170 27000 34260 27120
rect 34635 26310 34725 27090
rect 34635 25110 34725 26190
rect 35115 24510 35205 28290
rect 35355 27810 35445 27990
rect 35355 24510 35445 27690
rect 35595 27210 35685 29790
rect 36300 28695 36420 28710
rect 36555 28695 36645 30690
rect 36300 28605 36645 28695
rect 36300 28590 36420 28605
rect 36555 28110 36645 28605
rect 35595 26010 35685 27090
rect 35835 25410 35925 27390
rect 36555 26910 36645 27090
rect 36075 25110 36165 26490
rect 36555 25110 36645 26790
rect 34740 24405 35100 24495
rect 31275 20610 31365 21090
rect 29115 18705 29445 18795
rect 27915 15210 28005 16890
rect 28395 15810 28485 16290
rect 27915 10395 28005 12390
rect 28155 10710 28245 12990
rect 28395 11610 28485 15090
rect 28140 10590 28260 10710
rect 27915 10305 28245 10395
rect 25980 9120 26820 9210
rect 25890 8910 25980 9000
rect 26100 8910 26490 9000
rect 26730 9000 26820 9120
rect 26955 7710 27045 9090
rect 25950 6480 26040 7200
rect 26340 7200 26730 7290
rect 26970 7080 27060 7200
rect 26460 6990 27060 7080
rect 26970 6480 27060 6990
rect 27435 5910 27525 9090
rect 28155 7410 28245 10305
rect 28395 9810 28485 11490
rect 28395 7710 28485 8790
rect 28395 7110 28485 7590
rect 27675 6810 27765 6990
rect 27915 6510 28005 6690
rect 28635 2610 28725 15390
rect 29115 15210 29205 18705
rect 30795 18195 30885 19890
rect 32475 19110 32565 21690
rect 32715 21210 32805 21990
rect 33675 21810 33765 24090
rect 35115 21810 35205 23490
rect 31035 18510 31125 18990
rect 30795 18105 31125 18195
rect 31035 16710 31125 18105
rect 31020 16590 31140 16710
rect 31995 15810 32085 18690
rect 32715 18510 32805 21090
rect 32955 18510 33045 21090
rect 33435 19995 33525 20790
rect 33195 19905 33525 19995
rect 33195 19110 33285 19905
rect 33435 18810 33525 19590
rect 33675 18810 33765 21690
rect 34635 19410 34725 21090
rect 34875 18510 34965 20790
rect 35115 19710 35205 21690
rect 33675 17910 33765 18390
rect 30540 15210 30630 15720
rect 31290 15210 31380 15420
rect 30540 15120 31380 15210
rect 30315 13710 30405 15090
rect 30540 15000 30630 15120
rect 30870 14910 31260 15000
rect 31500 15000 31590 15720
rect 31380 14910 31470 15000
rect 31755 14010 31845 15090
rect 30300 13590 30420 13710
rect 29115 12810 29205 12990
rect 29355 10710 29445 12690
rect 30075 12210 30165 12390
rect 29340 10590 29460 10710
rect 31515 10110 31605 13290
rect 28875 8610 28965 9690
rect 29595 8910 29685 9090
rect 29595 6510 29685 8490
rect 30450 7200 30540 7290
rect 30330 6480 30420 7200
rect 30660 7200 31050 7290
rect 31290 7080 31380 7200
rect 30540 6990 31380 7080
rect 30540 6780 30630 6990
rect 31290 6480 31380 6990
rect 31515 6510 31605 9990
rect 31755 9210 31845 13890
rect 31995 13410 32085 15690
rect 32955 15210 33045 15990
rect 33675 15810 33765 17790
rect 35355 15510 35445 21090
rect 35595 20895 35685 24990
rect 35835 23910 35925 24690
rect 35595 20805 35925 20895
rect 35835 19110 35925 20805
rect 36075 20010 36165 24990
rect 36795 24510 36885 30690
rect 37275 27810 37365 33390
rect 37515 27810 37605 30090
rect 37755 28710 37845 30390
rect 37740 28590 37860 28710
rect 37995 28410 38085 33090
rect 38235 32910 38325 33090
rect 39675 31710 39765 32490
rect 39660 31590 39780 31710
rect 38235 30510 38325 30990
rect 38475 29910 38565 30990
rect 36555 23910 36645 24390
rect 35595 18810 35685 18990
rect 35835 17010 35925 18990
rect 36315 18510 36405 22290
rect 36555 21810 36645 23790
rect 37035 22410 37125 27690
rect 38475 27510 38565 29790
rect 39435 27810 39525 31590
rect 40155 30195 40245 33390
rect 41115 33210 41205 37290
rect 41355 33510 41445 36090
rect 42075 34110 42165 36990
rect 42315 36210 42405 36390
rect 41595 33810 41685 33990
rect 41355 33210 41445 33390
rect 42075 33210 42165 33690
rect 43515 33210 43605 41790
rect 43755 39210 43845 39690
rect 43995 39210 44085 42390
rect 44715 38910 44805 42990
rect 44955 42210 45045 42390
rect 43755 37410 43845 38490
rect 43755 37110 43845 37290
rect 43995 37110 44085 37290
rect 44715 36810 44805 36990
rect 44955 34710 45045 42090
rect 45195 39810 45285 43005
rect 45675 41610 45765 43305
rect 46050 43200 46140 43290
rect 45930 42480 46020 43200
rect 46260 43200 46650 43290
rect 46890 43080 46980 43200
rect 47730 43200 47820 43290
rect 46140 42990 46980 43080
rect 46140 42780 46230 42990
rect 46890 42480 46980 42990
rect 46155 39210 46245 42390
rect 46635 39510 46725 42090
rect 46875 39810 46965 41490
rect 46875 39210 46965 39690
rect 47115 39210 47205 42990
rect 47355 42510 47445 42990
rect 47610 42480 47700 43200
rect 47940 43200 48330 43290
rect 48570 43080 48660 43200
rect 47820 42990 48660 43080
rect 47820 42780 47910 42990
rect 48570 42480 48660 42990
rect 48795 41910 48885 42990
rect 45195 37710 45285 39090
rect 45180 37590 45300 37710
rect 46635 36510 46725 37290
rect 44940 34590 45060 34710
rect 43995 32010 44085 33090
rect 44490 33000 44580 33720
rect 44700 33210 44790 33420
rect 45450 33210 45540 33720
rect 46635 33510 46725 36390
rect 46875 35010 46965 39090
rect 47835 38910 47925 39390
rect 49755 38910 49845 39090
rect 51270 38160 52260 44040
rect 51270 38040 51330 38160
rect 52200 38040 52260 38160
rect 47595 36510 47685 36990
rect 49755 36810 49845 36990
rect 47595 33510 47685 33690
rect 48075 33510 48165 33690
rect 44700 33120 45540 33210
rect 44610 32910 44700 33000
rect 44820 32910 45210 33000
rect 45450 33000 45540 33120
rect 41355 31410 41445 31890
rect 43275 31110 43365 31290
rect 43995 31110 44085 31290
rect 40875 30510 40965 30990
rect 41595 30510 41685 30690
rect 40155 30105 40485 30195
rect 40395 28710 40485 30105
rect 40380 28590 40500 28710
rect 42075 27810 42165 27990
rect 38715 26910 38805 27090
rect 39195 25710 39285 27090
rect 39435 25695 39525 27690
rect 39930 27000 40020 27720
rect 40140 27210 40230 27420
rect 40890 27210 40980 27720
rect 42795 27210 42885 30990
rect 43515 30810 43605 30990
rect 43755 30810 43845 30990
rect 43755 30210 43845 30690
rect 43995 29910 44085 30690
rect 43515 27210 43605 27390
rect 43755 27210 43845 27990
rect 40140 27120 40980 27210
rect 40050 26910 40140 27000
rect 40260 26910 40650 27000
rect 40890 27000 40980 27120
rect 39435 25605 39765 25695
rect 39195 25410 39285 25590
rect 39435 23910 39525 24390
rect 39675 24210 39765 25605
rect 41115 25410 41205 27090
rect 43515 26610 43605 27090
rect 42555 25410 42645 25590
rect 43995 25410 44085 29790
rect 44475 27210 44565 31890
rect 45675 31710 45765 33090
rect 45915 32910 46005 33390
rect 46155 33210 46245 33390
rect 48315 33210 48405 36390
rect 49755 36195 49845 36690
rect 49515 36105 49845 36195
rect 49515 33210 49605 36105
rect 50475 35310 50565 36540
rect 48075 32910 48165 33090
rect 44715 25710 44805 27390
rect 44955 27210 45045 30390
rect 45195 27810 45285 31290
rect 46635 31110 46725 31290
rect 48450 31200 48540 31290
rect 46155 30510 46245 30690
rect 45915 25710 46005 27090
rect 46155 25410 46245 27390
rect 46635 26895 46725 27690
rect 47355 27510 47445 30990
rect 48330 30480 48420 31200
rect 48660 31200 49050 31290
rect 49290 31080 49380 31200
rect 48540 30990 49380 31080
rect 48540 30780 48630 30990
rect 49290 30480 49380 30990
rect 49515 30810 49605 33090
rect 47595 28710 47685 30090
rect 47580 28590 47700 28710
rect 49140 27705 49365 27795
rect 46635 26805 46860 26895
rect 43755 24810 43845 25290
rect 36555 19710 36645 21690
rect 37050 21000 37140 21720
rect 37260 21210 37350 21420
rect 38010 21210 38100 21720
rect 39675 21495 39765 24090
rect 39675 21405 40005 21495
rect 37260 21120 38100 21210
rect 37170 20910 37260 21000
rect 37380 20910 37770 21000
rect 38010 21000 38100 21120
rect 37275 19110 37365 19590
rect 36315 15810 36405 18390
rect 36795 18210 36885 18390
rect 36780 18090 36900 18210
rect 37275 17610 37365 18990
rect 37515 18810 37605 19890
rect 39675 19410 39765 21090
rect 34635 15210 34725 15390
rect 33300 15105 33660 15195
rect 33195 14910 33285 15090
rect 35595 14910 35685 15690
rect 32235 9210 32325 12090
rect 32475 9810 32565 12990
rect 32475 9210 32565 9690
rect 32715 7710 32805 14790
rect 34395 14310 34485 14790
rect 35835 14610 35925 14790
rect 33330 13200 33420 13290
rect 33210 12480 33300 13200
rect 33540 13200 33930 13290
rect 34170 13080 34260 13200
rect 34635 13110 34725 13290
rect 33420 12990 34260 13080
rect 33420 12780 33510 12990
rect 34170 12480 34260 12990
rect 33660 11490 33780 11610
rect 33675 9810 33765 11490
rect 35595 11295 35685 12990
rect 36315 11910 36405 14790
rect 36780 14490 36900 14610
rect 36555 13110 36645 13290
rect 36795 13110 36885 14490
rect 35355 11205 35685 11295
rect 33195 9210 33285 9690
rect 33420 9210 33510 9720
rect 33420 9120 34020 9210
rect 33420 9000 33510 9120
rect 33750 8910 34140 9000
rect 34440 9000 34530 9720
rect 35355 9210 35445 11205
rect 33900 8490 34020 8610
rect 33915 7995 34005 8490
rect 33675 7905 34005 7995
rect 30555 0 30645 6390
rect 32475 6210 32565 6990
rect 33675 6810 33765 7905
rect 35115 7110 35205 7290
rect 35355 7110 35445 7590
rect 33675 6510 33765 6690
rect 35595 2910 35685 9990
rect 36315 9210 36405 11790
rect 37035 10710 37125 12990
rect 37515 12510 37605 18690
rect 37755 15810 37845 18090
rect 37995 16710 38085 18990
rect 37980 16590 38100 16710
rect 37755 14910 37845 15090
rect 37995 13110 38085 15990
rect 38235 15510 38325 15690
rect 38235 15210 38325 15390
rect 38475 15210 38565 18390
rect 38955 18210 39045 18990
rect 39915 18510 40005 21405
rect 40395 20010 40485 21090
rect 40635 19410 40725 20790
rect 40395 18510 40485 18990
rect 40875 18510 40965 24390
rect 42315 24210 42405 24390
rect 42060 23490 42180 23610
rect 42075 21810 42165 23490
rect 46635 22710 46725 26490
rect 47355 25110 47445 27390
rect 48555 27210 48645 27390
rect 49275 27210 49365 27705
rect 49755 27210 49845 30990
rect 48555 25710 48645 27090
rect 49035 26910 49125 27090
rect 48540 25590 48660 25710
rect 48210 25200 48300 25290
rect 47835 23610 47925 24990
rect 48090 24480 48180 25200
rect 48420 25200 48810 25290
rect 49050 25080 49140 25200
rect 48300 24990 49140 25080
rect 48300 24780 48390 24990
rect 49050 24480 49140 24990
rect 46620 22590 46740 22710
rect 41115 19410 41205 21690
rect 42315 20910 42405 21090
rect 41580 20490 41700 20610
rect 41595 19710 41685 20490
rect 43515 19995 43605 21090
rect 43755 20910 43845 21090
rect 43515 19905 43845 19995
rect 42075 19110 42165 19590
rect 42315 18810 42405 19890
rect 43755 18810 43845 19905
rect 43995 19110 44085 21690
rect 44490 21000 44580 21720
rect 44700 21210 44790 21420
rect 45450 21210 45540 21720
rect 46140 21210 46230 21720
rect 46890 21210 46980 21420
rect 44700 21120 45540 21210
rect 44610 20910 44700 21000
rect 44820 20910 45210 21000
rect 45450 21000 45540 21120
rect 46140 21120 46980 21210
rect 44955 19995 45045 20490
rect 44715 19905 45045 19995
rect 44715 19110 44805 19905
rect 44475 18810 44565 18990
rect 44715 18810 44805 18990
rect 39435 16110 39525 18390
rect 40875 17910 40965 18390
rect 38715 13110 38805 15390
rect 38940 15210 39030 15720
rect 39690 15210 39780 15420
rect 38940 15120 39780 15210
rect 38940 15000 39030 15120
rect 39270 14910 39660 15000
rect 39900 15000 39990 15720
rect 39780 14910 39870 15000
rect 39435 13110 39525 14490
rect 40875 13695 40965 17790
rect 42315 15810 42405 18690
rect 41355 15210 41445 15390
rect 41595 14910 41685 15090
rect 41850 15000 41940 15720
rect 42060 15210 42150 15420
rect 42810 15210 42900 15720
rect 42060 15120 42900 15210
rect 41970 14910 42060 15000
rect 42180 14910 42570 15000
rect 42810 15000 42900 15120
rect 40875 13605 41205 13695
rect 41115 13110 41205 13605
rect 37995 12510 38085 12690
rect 37020 10590 37140 10710
rect 37275 9810 37365 9990
rect 37515 9810 37605 12390
rect 37995 11595 38085 12390
rect 37755 11505 38085 11595
rect 37755 10710 37845 11505
rect 37740 10590 37860 10710
rect 36795 9495 36885 9690
rect 36795 9405 37125 9495
rect 36555 6510 36645 7590
rect 36795 7410 36885 7590
rect 37035 6210 37125 9405
rect 38475 9210 38565 12990
rect 38715 12810 38805 12990
rect 38475 7710 38565 9090
rect 38715 7110 38805 12690
rect 39435 12510 39525 12990
rect 39435 9495 39525 12390
rect 39915 9510 40005 12990
rect 41595 12210 41685 12990
rect 39435 9405 39765 9495
rect 38955 7110 39045 9090
rect 39675 7110 39765 9405
rect 39915 9210 40005 9390
rect 40875 7710 40965 9690
rect 41115 9210 41205 9990
rect 39435 6810 39525 6990
rect 36555 0 36645 6090
rect 40395 300 40485 7590
rect 40875 7110 40965 7590
rect 42075 7110 42165 9690
rect 42555 9210 42645 14190
rect 43035 12210 43125 15090
rect 43275 14910 43365 18390
rect 43500 17490 43620 17610
rect 43515 15210 43605 17490
rect 43275 13110 43365 14790
rect 43755 12810 43845 15690
rect 43995 13110 44085 18690
rect 44475 15210 44565 15690
rect 44715 15210 44805 15390
rect 45195 15210 45285 20190
rect 45915 19710 46005 21090
rect 46140 21000 46230 21120
rect 46470 20910 46860 21000
rect 47100 21000 47190 21720
rect 47355 21210 47445 21390
rect 47835 21195 47925 23490
rect 47835 21105 48165 21195
rect 46980 20910 47070 21000
rect 46635 18810 46725 19890
rect 47355 19110 47445 21090
rect 47595 20010 47685 20790
rect 48075 19410 48165 21105
rect 49515 20295 49605 24990
rect 49275 20205 49605 20295
rect 48075 19110 48165 19290
rect 49275 18810 49365 20205
rect 49755 19710 49845 21090
rect 49995 20610 50085 21390
rect 49740 19590 49860 19710
rect 46635 18510 46725 18690
rect 48075 17895 48165 18690
rect 47835 17805 48165 17895
rect 46875 15810 46965 17490
rect 47835 16710 47925 17805
rect 47820 16590 47940 16710
rect 46635 13110 46725 15690
rect 43275 10710 43365 12690
rect 43755 11910 43845 12390
rect 43260 10590 43380 10710
rect 42555 8010 42645 9090
rect 42810 9000 42900 9720
rect 43020 9210 43110 9420
rect 43770 9210 43860 9720
rect 43995 9510 44085 12990
rect 44715 12510 44805 12690
rect 43020 9120 43860 9210
rect 42930 8910 43020 9000
rect 43140 8910 43530 9000
rect 43770 9000 43860 9120
rect 42555 7410 42645 7890
rect 40875 6510 40965 6990
rect 40380 210 40485 300
rect 40380 0 40470 210
rect 42555 0 42645 6990
rect 43995 6810 44085 9090
rect 44235 6810 44325 6990
rect 44475 6810 44565 9390
rect 45195 9210 45285 12990
rect 45450 9000 45540 9720
rect 45660 9210 45750 9420
rect 46410 9210 46500 9720
rect 45660 9120 46500 9210
rect 45570 8910 45660 9000
rect 45780 8910 46170 9000
rect 46410 9000 46500 9120
rect 46635 7410 46725 12390
rect 46875 9810 46965 15690
rect 48075 14910 48165 15090
rect 48315 13710 48405 13890
rect 48300 13590 48420 13710
rect 47595 9810 47685 12990
rect 47835 12510 47925 12690
rect 48795 12510 48885 15090
rect 49755 13110 49845 15390
rect 47595 9210 47685 9390
rect 48315 9210 48405 12390
rect 46875 6810 46965 9090
rect 43995 6510 44085 6690
rect 47355 6510 47445 7290
rect 48075 7110 48165 7890
rect 47835 6510 47925 6690
rect 48555 0 48645 12090
rect 49035 11895 49125 12390
rect 49035 11805 49365 11895
rect 49275 10710 49365 11805
rect 49755 11295 49845 12990
rect 49995 12810 50085 15690
rect 50235 11610 50325 12540
rect 49515 11205 49845 11295
rect 49260 10590 49380 10710
rect 49515 9210 49605 11205
rect 50955 5310 51045 32490
rect 51270 32160 52260 38040
rect 51270 32040 51330 32160
rect 52200 32040 52260 32160
rect 51270 26160 52260 32040
rect 51270 26040 51330 26160
rect 52200 26040 52260 26160
rect 51270 20160 52260 26040
rect 51270 20040 51330 20160
rect 52200 20040 52260 20160
rect 51270 14160 52260 20040
rect 51270 14040 51330 14160
rect 52200 14040 52260 14160
rect 51270 8160 52260 14040
rect 51270 8040 51330 8160
rect 52200 8040 52260 8160
rect 51270 3976 52260 8040
rect 51270 3104 51330 3976
rect 52200 3104 52260 3976
rect 51270 3045 52260 3104
rect 53250 41160 54240 47204
rect 54450 42810 54540 49200
rect 53250 41040 53310 41160
rect 54180 41040 54240 41160
rect 53250 35160 54240 41040
rect 53250 35040 53310 35160
rect 54180 35040 54240 35160
rect 53250 29160 54240 35040
rect 53250 29040 53310 29160
rect 54180 29040 54240 29160
rect 53250 23160 54240 29040
rect 53250 23040 53310 23160
rect 54180 23040 54240 23160
rect 53250 17160 54240 23040
rect 53250 17040 53310 17160
rect 54180 17040 54240 17160
rect 53250 11160 54240 17040
rect 53250 11040 53310 11160
rect 54180 11040 54240 11160
rect 53250 5160 54240 11040
rect 53250 5040 53310 5160
rect 54180 5040 54240 5160
rect 53250 1996 54240 5040
rect 53250 1124 53310 1996
rect 54180 1124 54240 1996
rect 54555 1140 54645 11790
rect 53250 1065 54240 1124
<< m3contact >>
rect 2460 38790 2580 38910
rect 780 26190 900 26310
rect 9420 43890 9540 44010
rect 7500 43590 7620 43710
rect 6540 42990 6660 43110
rect 7260 42990 7380 43110
rect 8700 42990 8820 43110
rect 6780 42690 6900 42810
rect 5580 42390 5700 42510
rect 6540 42390 6660 42510
rect 7740 42390 7860 42510
rect 8460 42390 8580 42510
rect 8940 42390 9060 42510
rect 12300 43290 12420 43410
rect 13020 43290 13140 43410
rect 10380 42990 10500 43110
rect 10860 42990 10980 43110
rect 11340 42990 11460 43110
rect 9660 42690 9780 42810
rect 9660 42390 9780 42510
rect 9660 39390 9780 39510
rect 5340 38040 5460 38160
rect 2700 37590 2820 37710
rect 2700 37290 2820 37410
rect 2460 15990 2580 16110
rect 2700 13290 2820 13410
rect 2700 6390 2820 6510
rect 6060 39090 6180 39210
rect 7500 39090 7620 39210
rect 6780 36990 6900 37110
rect 7260 36990 7380 37110
rect 5580 36390 5700 36510
rect 7020 36390 7140 36510
rect 7260 33690 7380 33810
rect 6540 32640 6660 32760
rect 8220 36390 8340 36510
rect 9180 36390 9300 36510
rect 11340 39990 11460 40110
rect 13740 42990 13860 43110
rect 13980 42690 14100 42810
rect 12780 39990 12900 40110
rect 13020 39390 13140 39510
rect 13260 39090 13380 39210
rect 12300 37590 12420 37710
rect 10860 37290 10980 37410
rect 12060 37290 12180 37410
rect 10860 36990 10980 37110
rect 10860 36690 10980 36810
rect 11340 36690 11460 36810
rect 13020 36990 13140 37110
rect 7740 33690 7860 33810
rect 6060 31590 6180 31710
rect 7020 31590 7140 31710
rect 6300 31290 6420 31410
rect 5340 30390 5460 30510
rect 6060 27240 6180 27360
rect 10140 36090 10260 36210
rect 12780 33990 12900 34110
rect 8220 31290 8340 31410
rect 7980 30990 8100 31110
rect 9180 30990 9300 31110
rect 8220 30690 8340 30810
rect 8460 30390 8580 30510
rect 7740 27390 7860 27510
rect 11580 32790 11700 32910
rect 10860 32190 10980 32310
rect 11820 32190 11940 32310
rect 9660 30990 9780 31110
rect 10140 30690 10260 30810
rect 9420 30090 9540 30210
rect 9180 29490 9300 29610
rect 9900 29490 10020 29610
rect 8700 27390 8820 27510
rect 9180 27390 9300 27510
rect 8700 26790 8820 26910
rect 11820 30390 11940 30510
rect 11340 27690 11460 27810
rect 12060 30090 12180 30210
rect 12060 29790 12180 29910
rect 12540 27990 12660 28110
rect 18060 46890 18180 47010
rect 15180 46590 15300 46710
rect 14700 42990 14820 43110
rect 14460 39990 14580 40110
rect 14220 39090 14340 39210
rect 13500 33090 13620 33210
rect 13980 33090 14100 33210
rect 13740 30690 13860 30810
rect 13020 30390 13140 30510
rect 17100 43290 17220 43410
rect 15900 42690 16020 42810
rect 17340 42690 17460 42810
rect 15900 42390 16020 42510
rect 15660 41190 15780 41310
rect 14700 36990 14820 37110
rect 14940 36390 15060 36510
rect 16140 38490 16260 38610
rect 15420 36990 15540 37110
rect 15180 34290 15300 34410
rect 15180 33090 15300 33210
rect 17580 38790 17700 38910
rect 17100 37290 17220 37410
rect 16380 36990 16500 37110
rect 16140 36390 16260 36510
rect 16140 36090 16260 36210
rect 16860 33390 16980 33510
rect 15900 33090 16020 33210
rect 16620 33090 16740 33210
rect 15660 32790 15780 32910
rect 16380 32490 16500 32610
rect 12780 27690 12900 27810
rect 13260 27690 13380 27810
rect 15180 27690 15300 27810
rect 17340 33690 17460 33810
rect 22380 43890 22500 44010
rect 18540 43590 18660 43710
rect 19020 43290 19140 43410
rect 18060 42390 18180 42510
rect 18300 39090 18420 39210
rect 18780 39090 18900 39210
rect 20220 43290 20340 43410
rect 19260 42390 19380 42510
rect 19740 42390 19860 42510
rect 20700 42690 20820 42810
rect 19500 39390 19620 39510
rect 23340 43590 23460 43710
rect 27660 43590 27780 43710
rect 28620 43590 28740 43710
rect 31500 43290 31620 43410
rect 28140 42990 28260 43110
rect 28860 42990 28980 43110
rect 32220 42990 32340 43110
rect 25020 42390 25140 42510
rect 25980 42390 26100 42510
rect 25740 42090 25860 42210
rect 22620 40890 22740 41010
rect 24060 40890 24180 41010
rect 21420 39390 21540 39510
rect 20940 39090 21060 39210
rect 18540 36990 18660 37110
rect 18780 34290 18900 34410
rect 18540 33690 18660 33810
rect 17580 33390 17700 33510
rect 17100 32490 17220 32610
rect 16860 31590 16980 31710
rect 17340 31590 17460 31710
rect 17100 30090 17220 30210
rect 17580 30090 17700 30210
rect 15900 27690 16020 27810
rect 13260 27390 13380 27510
rect 15420 27390 15540 27510
rect 11100 27090 11220 27210
rect 12540 27090 12660 27210
rect 10380 26790 10500 26910
rect 7740 26490 7860 26610
rect 9420 25890 9540 26010
rect 10140 25890 10260 26010
rect 5340 24990 5460 25110
rect 8460 25290 8580 25410
rect 9420 25290 9540 25410
rect 7020 24990 7140 25110
rect 8700 24990 8820 25110
rect 6780 24690 6900 24810
rect 6060 21990 6180 22110
rect 5340 21090 5460 21210
rect 7500 24390 7620 24510
rect 8700 24390 8820 24510
rect 12060 25290 12180 25410
rect 13020 25290 13140 25410
rect 10860 24990 10980 25110
rect 10140 24690 10260 24810
rect 12060 23490 12180 23610
rect 9660 21690 9780 21810
rect 10380 21690 10500 21810
rect 7020 21390 7140 21510
rect 10380 21390 10500 21510
rect 7020 21090 7140 21210
rect 10140 21090 10260 21210
rect 6780 20790 6900 20910
rect 9660 20790 9780 20910
rect 8940 20490 9060 20610
rect 11820 21090 11940 21210
rect 11580 20490 11700 20610
rect 10860 17490 10980 17610
rect 8460 16590 8580 16710
rect 9420 16290 9540 16410
rect 6780 15690 6900 15810
rect 6060 15090 6180 15210
rect 7020 13590 7140 13710
rect 5340 11040 5460 11160
rect 6300 9990 6420 10110
rect 5580 9690 5700 9810
rect 6540 9690 6660 9810
rect 6780 9390 6900 9510
rect 5580 6990 5700 7110
rect 9420 15690 9540 15810
rect 9180 15390 9300 15510
rect 10140 15390 10260 15510
rect 10860 15090 10980 15210
rect 9660 14490 9780 14610
rect 8220 12990 8340 13110
rect 9420 12990 9540 13110
rect 16620 27090 16740 27210
rect 15180 26490 15300 26610
rect 15420 26190 15540 26310
rect 17820 29490 17940 29610
rect 20940 36990 21060 37110
rect 21420 36990 21540 37110
rect 19500 36690 19620 36810
rect 19980 36390 20100 36510
rect 21420 36390 21540 36510
rect 19740 33990 19860 34110
rect 21420 36090 21540 36210
rect 21180 33690 21300 33810
rect 19020 33090 19140 33210
rect 19500 32790 19620 32910
rect 21180 32790 21300 32910
rect 30540 42690 30660 42810
rect 31260 42690 31380 42810
rect 31980 42690 32100 42810
rect 32460 42690 32580 42810
rect 27900 42390 28020 42510
rect 29580 42390 29700 42510
rect 27180 42090 27300 42210
rect 28860 41190 28980 41310
rect 26220 40590 26340 40710
rect 24060 39390 24180 39510
rect 21900 38790 22020 38910
rect 23820 39090 23940 39210
rect 24300 39090 24420 39210
rect 27180 39390 27300 39510
rect 27180 39090 27300 39210
rect 23580 38790 23700 38910
rect 24780 38790 24900 38910
rect 25740 38790 25860 38910
rect 22380 37290 22500 37410
rect 24300 37290 24420 37410
rect 23820 36990 23940 37110
rect 23100 36090 23220 36210
rect 22860 35790 22980 35910
rect 21660 32190 21780 32310
rect 19260 31290 19380 31410
rect 19020 30690 19140 30810
rect 21180 31290 21300 31410
rect 22860 31290 22980 31410
rect 20940 30990 21060 31110
rect 21660 30990 21780 31110
rect 22620 30990 22740 31110
rect 19980 30690 20100 30810
rect 21180 30390 21300 30510
rect 21900 30390 22020 30510
rect 20940 30090 21060 30210
rect 19740 29490 19860 29610
rect 17820 27690 17940 27810
rect 19260 27390 19380 27510
rect 18060 27090 18180 27210
rect 17100 25890 17220 26010
rect 17580 25890 17700 26010
rect 13500 24990 13620 25110
rect 14220 24990 14340 25110
rect 15420 24990 15540 25110
rect 13500 24690 13620 24810
rect 13980 23490 14100 23610
rect 15660 24690 15780 24810
rect 14220 22590 14340 22710
rect 11580 18390 11700 18510
rect 15660 20190 15780 20310
rect 13260 19290 13380 19410
rect 12540 15990 12660 16110
rect 11580 14790 11700 14910
rect 13020 15690 13140 15810
rect 12540 14790 12660 14910
rect 11820 14490 11940 14610
rect 11100 14190 11220 14310
rect 11580 14190 11700 14310
rect 12780 14190 12900 14310
rect 9900 13290 10020 13410
rect 10860 12990 10980 13110
rect 12780 12990 12900 13110
rect 7260 9990 7380 10110
rect 8460 9990 8580 10110
rect 7740 9090 7860 9210
rect 8460 9390 8580 9510
rect 9420 9390 9540 9510
rect 11340 12390 11460 12510
rect 12540 12390 12660 12510
rect 12540 9690 12660 9810
rect 9900 9390 10020 9510
rect 10380 9390 10500 9510
rect 9660 9090 9780 9210
rect 10140 9090 10260 9210
rect 8220 7290 8340 7410
rect 10140 7290 10260 7410
rect 10380 6990 10500 7110
rect 12300 6990 12420 7110
rect 12780 6990 12900 7110
rect 6540 6090 6660 6210
rect 7020 6090 7140 6210
rect 7740 6090 7860 6210
rect 6300 720 6420 840
rect 9900 6690 10020 6810
rect 9420 6390 9540 6510
rect 10380 6390 10500 6510
rect 10860 6390 10980 6510
rect 11820 6390 11940 6510
rect 12300 6390 12420 6510
rect 12780 6390 12900 6510
rect 13500 18690 13620 18810
rect 14940 19290 15060 19410
rect 15420 18990 15540 19110
rect 15660 18690 15780 18810
rect 16140 17490 16260 17610
rect 13980 16290 14100 16410
rect 16380 15990 16500 16110
rect 14220 15690 14340 15810
rect 14940 15690 15060 15810
rect 14700 15390 14820 15510
rect 13740 14790 13860 14910
rect 15660 15390 15780 15510
rect 16860 15690 16980 15810
rect 16620 15090 16740 15210
rect 18780 26790 18900 26910
rect 18060 22890 18180 23010
rect 18060 22290 18180 22410
rect 22140 29790 22260 29910
rect 25020 36990 25140 37110
rect 25740 36990 25860 37110
rect 28140 38790 28260 38910
rect 27900 36990 28020 37110
rect 28380 36990 28500 37110
rect 24780 34290 24900 34410
rect 26220 36390 26340 36510
rect 27180 36390 27300 36510
rect 24540 33690 24660 33810
rect 25260 33690 25380 33810
rect 21660 27990 21780 28110
rect 23100 27990 23220 28110
rect 21660 27690 21780 27810
rect 23820 33090 23940 33210
rect 24060 30990 24180 31110
rect 23580 27990 23700 28110
rect 24060 27690 24180 27810
rect 24780 33090 24900 33210
rect 25260 32790 25380 32910
rect 25740 33090 25860 33210
rect 26700 33390 26820 33510
rect 31500 42390 31620 42510
rect 32220 42390 32340 42510
rect 31260 42090 31380 42210
rect 36540 43590 36660 43710
rect 40140 43590 40260 43710
rect 45660 43590 45780 43710
rect 46380 43590 46500 43710
rect 34620 42990 34740 43110
rect 35100 42990 35220 43110
rect 33660 42690 33780 42810
rect 33180 42090 33300 42210
rect 30780 38490 30900 38610
rect 31260 37590 31380 37710
rect 32940 37590 33060 37710
rect 30060 37290 30180 37410
rect 31020 37290 31140 37410
rect 32700 37290 32820 37410
rect 28380 36090 28500 36210
rect 28860 36090 28980 36210
rect 28380 35190 28500 35310
rect 29580 35790 29700 35910
rect 30540 33990 30660 34110
rect 32940 36990 33060 37110
rect 31980 36690 32100 36810
rect 32460 36690 32580 36810
rect 31260 36390 31380 36510
rect 31740 36390 31860 36510
rect 31740 33690 31860 33810
rect 32700 33990 32820 34110
rect 32700 33690 32820 33810
rect 31020 33390 31140 33510
rect 31740 33390 31860 33510
rect 34140 40590 34260 40710
rect 33420 39090 33540 39210
rect 33420 38790 33540 38910
rect 35100 39090 35220 39210
rect 35580 39090 35700 39210
rect 33180 36390 33300 36510
rect 35100 36990 35220 37110
rect 33660 36390 33780 36510
rect 34380 36390 34500 36510
rect 33420 34290 33540 34410
rect 33180 33090 33300 33210
rect 29100 32790 29220 32910
rect 26220 32190 26340 32310
rect 25500 31290 25620 31410
rect 25980 30990 26100 31110
rect 25740 30690 25860 30810
rect 25500 29490 25620 29610
rect 25500 27990 25620 28110
rect 23340 27390 23460 27510
rect 24540 27390 24660 27510
rect 25500 27390 25620 27510
rect 20700 27090 20820 27210
rect 21180 27090 21300 27210
rect 25260 27090 25380 27210
rect 22380 24990 22500 25110
rect 18540 22890 18660 23010
rect 17580 21090 17700 21210
rect 18300 21090 18420 21210
rect 17340 18390 17460 18510
rect 16620 14490 16740 14610
rect 17100 14490 17220 14610
rect 17820 14790 17940 14910
rect 16860 13890 16980 14010
rect 17580 13890 17700 14010
rect 15900 13290 16020 13410
rect 15180 12390 15300 12510
rect 15180 10590 15300 10710
rect 16380 9390 16500 9510
rect 16380 9090 16500 9210
rect 19740 23490 19860 23610
rect 20220 22890 20340 23010
rect 21180 22890 21300 23010
rect 19740 22290 19860 22410
rect 18540 20790 18660 20910
rect 21180 22590 21300 22710
rect 20220 20790 20340 20910
rect 19500 20490 19620 20610
rect 19740 20190 19860 20310
rect 18540 18990 18660 19110
rect 18300 18690 18420 18810
rect 22140 21390 22260 21510
rect 24060 26490 24180 26610
rect 25740 26490 25860 26610
rect 25500 25890 25620 26010
rect 23100 24390 23220 24510
rect 23580 24390 23700 24510
rect 22620 21690 22740 21810
rect 23100 21390 23220 21510
rect 20460 20490 20580 20610
rect 20940 18690 21060 18810
rect 20940 18390 21060 18510
rect 21420 18390 21540 18510
rect 19500 17790 19620 17910
rect 18300 17490 18420 17610
rect 18540 15690 18660 15810
rect 18780 15090 18900 15210
rect 18060 13590 18180 13710
rect 17100 12990 17220 13110
rect 14220 6690 14340 6810
rect 15900 6990 16020 7110
rect 13260 6390 13380 6510
rect 15420 6390 15540 6510
rect 13020 6090 13140 6210
rect 8460 5640 8580 5760
rect 19020 12990 19140 13110
rect 19020 12690 19140 12810
rect 18060 10590 18180 10710
rect 18780 9990 18900 10110
rect 17340 9090 17460 9210
rect 19500 14190 19620 14310
rect 20460 15990 20580 16110
rect 21420 15690 21540 15810
rect 20220 15090 20340 15210
rect 20220 13590 20340 13710
rect 20220 13290 20340 13410
rect 19980 10890 20100 11010
rect 19260 9990 19380 10110
rect 19260 9090 19380 9210
rect 19020 8790 19140 8910
rect 22140 18990 22260 19110
rect 22620 18990 22740 19110
rect 22860 18690 22980 18810
rect 23580 16890 23700 17010
rect 22140 15690 22260 15810
rect 22620 15390 22740 15510
rect 21900 14790 22020 14910
rect 23580 15090 23700 15210
rect 22380 13290 22500 13410
rect 21660 12690 21780 12810
rect 21420 12390 21540 12510
rect 22620 12390 22740 12510
rect 20940 10890 21060 11010
rect 21900 9390 22020 9510
rect 20940 9090 21060 9210
rect 21660 9090 21780 9210
rect 20940 8790 21060 8910
rect 23340 9690 23460 9810
rect 24300 24990 24420 25110
rect 24540 23790 24660 23910
rect 24060 19890 24180 20010
rect 33660 33690 33780 33810
rect 35100 36090 35220 36210
rect 34860 34590 34980 34710
rect 35340 35790 35460 35910
rect 35100 33990 35220 34110
rect 26940 31290 27060 31410
rect 27420 31290 27540 31410
rect 29820 31290 29940 31410
rect 26700 30390 26820 30510
rect 27180 30690 27300 30810
rect 26940 29190 27060 29310
rect 27420 30390 27540 30510
rect 29100 30990 29220 31110
rect 32220 31290 32340 31410
rect 29100 30690 29220 30810
rect 29580 30690 29700 30810
rect 28620 30390 28740 30510
rect 28620 30090 28740 30210
rect 28380 29790 28500 29910
rect 27660 29490 27780 29610
rect 27180 24690 27300 24810
rect 25500 23490 25620 23610
rect 25500 21690 25620 21810
rect 26220 21390 26340 21510
rect 26700 21390 26820 21510
rect 24540 19890 24660 20010
rect 25980 19890 26100 20010
rect 24540 19590 24660 19710
rect 26940 19590 27060 19710
rect 24300 18990 24420 19110
rect 24300 16890 24420 17010
rect 24060 16590 24180 16710
rect 24060 15390 24180 15510
rect 26220 19290 26340 19410
rect 27180 19290 27300 19410
rect 26220 18990 26340 19110
rect 25260 17490 25380 17610
rect 26460 18690 26580 18810
rect 26940 18690 27060 18810
rect 27420 18090 27540 18210
rect 24780 16590 24900 16710
rect 25980 16590 26100 16710
rect 26460 16590 26580 16710
rect 24540 15990 24660 16110
rect 25260 15990 25380 16110
rect 24300 11790 24420 11910
rect 25020 15690 25140 15810
rect 25500 15390 25620 15510
rect 27180 15090 27300 15210
rect 26700 13290 26820 13410
rect 24780 12990 24900 13110
rect 26220 12990 26340 13110
rect 26700 12990 26820 13110
rect 24780 11790 24900 11910
rect 24060 9090 24180 9210
rect 23820 8790 23940 8910
rect 18780 8490 18900 8610
rect 17820 7590 17940 7710
rect 18540 7590 18660 7710
rect 21180 8490 21300 8610
rect 18540 6090 18660 6210
rect 20700 6090 20820 6210
rect 18540 5190 18660 5310
rect 24540 8790 24660 8910
rect 24300 6990 24420 7110
rect 23340 5790 23460 5910
rect 12540 750 12660 870
rect 25260 12690 25380 12810
rect 26940 12690 27060 12810
rect 25500 9690 25620 9810
rect 28380 27390 28500 27510
rect 30060 30090 30180 30210
rect 29100 29790 29220 29910
rect 28860 27390 28980 27510
rect 34620 32790 34740 32910
rect 33660 30390 33780 30510
rect 33900 29490 34020 29610
rect 33660 29190 33780 29310
rect 33180 27990 33300 28110
rect 32940 27690 33060 27810
rect 27900 24990 28020 25110
rect 30300 27390 30420 27510
rect 32220 27390 32340 27510
rect 31980 27090 32100 27210
rect 30780 26790 30900 26910
rect 30540 25290 30660 25410
rect 30540 24990 30660 25110
rect 29340 24690 29460 24810
rect 32460 26790 32580 26910
rect 31740 25290 31860 25410
rect 32700 25290 32820 25410
rect 29340 24390 29460 24510
rect 28140 23490 28260 23610
rect 29100 23490 29220 23610
rect 27900 21690 28020 21810
rect 28860 21690 28980 21810
rect 28860 21090 28980 21210
rect 30780 24090 30900 24210
rect 29820 21090 29940 21210
rect 30540 20490 30660 20610
rect 35100 33090 35220 33210
rect 35100 31590 35220 31710
rect 35100 31290 35220 31410
rect 35100 30390 35220 30510
rect 37260 42990 37380 43110
rect 38460 42990 38580 43110
rect 40860 43290 40980 43410
rect 41340 43290 41460 43410
rect 42540 43290 42660 43410
rect 36540 42690 36660 42810
rect 36060 39090 36180 39210
rect 35820 37590 35940 37710
rect 39180 39390 39300 39510
rect 38220 38790 38340 38910
rect 37500 38490 37620 38610
rect 37020 37290 37140 37410
rect 36300 36090 36420 36210
rect 36300 34890 36420 35010
rect 36300 33990 36420 34110
rect 35820 33090 35940 33210
rect 36540 33690 36660 33810
rect 37260 34590 37380 34710
rect 40860 39390 40980 39510
rect 41580 39390 41700 39510
rect 42300 39390 42420 39510
rect 38940 39090 39060 39210
rect 39900 39090 40020 39210
rect 44220 42990 44340 43110
rect 44700 42990 44820 43110
rect 44460 42690 44580 42810
rect 43500 41790 43620 41910
rect 40860 38790 40980 38910
rect 40620 38490 40740 38610
rect 39420 37590 39540 37710
rect 40380 37290 40500 37410
rect 39420 36390 39540 36510
rect 40380 35490 40500 35610
rect 37260 33390 37380 33510
rect 39420 33390 39540 33510
rect 40140 33390 40260 33510
rect 40860 33390 40980 33510
rect 37020 32490 37140 32610
rect 36780 30990 36900 31110
rect 36300 30690 36420 30810
rect 36780 30690 36900 30810
rect 36060 30390 36180 30510
rect 35100 30090 35220 30210
rect 35580 30090 35700 30210
rect 34860 29790 34980 29910
rect 35580 29790 35700 29910
rect 35100 28290 35220 28410
rect 34380 27090 34500 27210
rect 34620 26190 34740 26310
rect 33180 24990 33300 25110
rect 35340 27990 35460 28110
rect 36540 27990 36660 28110
rect 35820 27390 35940 27510
rect 35580 25890 35700 26010
rect 36060 27090 36180 27210
rect 36540 27090 36660 27210
rect 36540 26790 36660 26910
rect 36060 26490 36180 26610
rect 35580 24990 35700 25110
rect 33660 24390 33780 24510
rect 35340 24390 35460 24510
rect 31740 24090 31860 24210
rect 32940 24090 33060 24210
rect 33660 24090 33780 24210
rect 32700 21990 32820 22110
rect 31260 20490 31380 20610
rect 31020 20190 31140 20310
rect 30780 19890 30900 20010
rect 29580 18990 29700 19110
rect 28380 18390 28500 18510
rect 27900 16890 28020 17010
rect 27660 16290 27780 16410
rect 28380 16290 28500 16410
rect 28380 11490 28500 11610
rect 26460 7590 26580 7710
rect 26940 7590 27060 7710
rect 26220 7290 26340 7410
rect 28380 8790 28500 8910
rect 28380 7590 28500 7710
rect 27900 6990 28020 7110
rect 27660 6690 27780 6810
rect 27900 6390 28020 6510
rect 28380 6390 28500 6510
rect 27420 5790 27540 5910
rect 29340 18390 29460 18510
rect 35100 23490 35220 23610
rect 32700 21090 32820 21210
rect 31020 18990 31140 19110
rect 31980 18990 32100 19110
rect 31980 18690 32100 18810
rect 30060 15690 30180 15810
rect 33420 19590 33540 19710
rect 34620 19290 34740 19410
rect 33660 18690 33780 18810
rect 35100 19590 35220 19710
rect 32940 18390 33060 18510
rect 33660 18390 33780 18510
rect 33660 17790 33780 17910
rect 32940 15990 33060 16110
rect 31980 15690 32100 15810
rect 31740 13890 31860 14010
rect 31500 13290 31620 13410
rect 29580 12990 29700 13110
rect 29100 12690 29220 12810
rect 30780 12690 30900 12810
rect 30300 12390 30420 12510
rect 30060 12090 30180 12210
rect 31500 9990 31620 10110
rect 29580 9090 29700 9210
rect 31020 9090 31140 9210
rect 29100 8790 29220 8910
rect 29820 8790 29940 8910
rect 28860 8490 28980 8610
rect 29580 8490 29700 8610
rect 30060 6990 30180 7110
rect 30780 6690 30900 6810
rect 30540 6390 30660 6510
rect 35820 24690 35940 24810
rect 35820 23790 35940 23910
rect 39420 33090 39540 33210
rect 37740 30390 37860 30510
rect 38220 32790 38340 32910
rect 39900 32790 40020 32910
rect 39660 32490 39780 32610
rect 39420 31590 39540 31710
rect 38220 30990 38340 31110
rect 39180 30690 39300 30810
rect 38460 29790 38580 29910
rect 37980 28290 38100 28410
rect 36540 23790 36660 23910
rect 36300 23490 36420 23610
rect 36300 22290 36420 22410
rect 36060 19890 36180 20010
rect 36060 18990 36180 19110
rect 35580 18690 35700 18810
rect 39660 30690 39780 30810
rect 43260 36990 43380 37110
rect 41340 36090 41460 36210
rect 42300 36690 42420 36810
rect 42780 36690 42900 36810
rect 42300 36090 42420 36210
rect 43260 35490 43380 35610
rect 41580 33990 41700 34110
rect 42060 33990 42180 34110
rect 41820 33690 41940 33810
rect 41340 33390 41460 33510
rect 42300 33390 42420 33510
rect 43740 39090 43860 39210
rect 44940 42690 45060 42810
rect 44940 42090 45060 42210
rect 43740 38490 43860 38610
rect 43980 37290 44100 37410
rect 43740 36990 43860 37110
rect 44700 36990 44820 37110
rect 45420 42990 45540 43110
rect 46140 42390 46260 42510
rect 45660 41490 45780 41610
rect 45900 39390 46020 39510
rect 46620 42090 46740 42210
rect 46860 41490 46980 41610
rect 46860 39690 46980 39810
rect 46380 39390 46500 39510
rect 47340 42390 47460 42510
rect 48780 41790 48900 41910
rect 49260 39690 49380 39810
rect 45180 39090 45300 39210
rect 47100 39090 47220 39210
rect 45420 38490 45540 38610
rect 46620 37290 46740 37410
rect 45420 36990 45540 37110
rect 43740 33690 43860 33810
rect 41100 33090 41220 33210
rect 42060 33090 42180 33210
rect 43980 33090 44100 33210
rect 41340 32490 41460 32610
rect 48060 39090 48180 39210
rect 47820 38790 47940 38910
rect 49740 38790 49860 38910
rect 48060 36990 48180 37110
rect 47820 36690 47940 36810
rect 49740 36690 49860 36810
rect 47580 36390 47700 36510
rect 48300 36390 48420 36510
rect 49260 36390 49380 36510
rect 46860 34890 46980 35010
rect 47340 33690 47460 33810
rect 48060 33690 48180 33810
rect 46140 33390 46260 33510
rect 46620 33390 46740 33510
rect 47580 33390 47700 33510
rect 41340 31890 41460 32010
rect 43980 31890 44100 32010
rect 44460 31890 44580 32010
rect 43260 31290 43380 31410
rect 43980 31290 44100 31410
rect 40860 30990 40980 31110
rect 42780 30990 42900 31110
rect 43500 30990 43620 31110
rect 41580 30690 41700 30810
rect 40380 30390 40500 30510
rect 42060 27990 42180 28110
rect 38940 27690 39060 27810
rect 38460 27390 38580 27510
rect 38460 27090 38580 27210
rect 38700 26790 38820 26910
rect 39180 25590 39300 25710
rect 43740 30690 43860 30810
rect 43740 30090 43860 30210
rect 43980 29790 44100 29910
rect 43740 27990 43860 28110
rect 41340 27090 41460 27210
rect 43500 27090 43620 27210
rect 38700 25290 38820 25410
rect 39180 25290 39300 25410
rect 38940 24990 39060 25110
rect 39420 24990 39540 25110
rect 37980 24390 38100 24510
rect 43500 26490 43620 26610
rect 42540 25590 42660 25710
rect 50460 36540 50580 36660
rect 50460 35190 50580 35310
rect 46620 33090 46740 33210
rect 45900 32790 46020 32910
rect 48060 32790 48180 32910
rect 45180 31290 45300 31410
rect 46620 31290 46740 31410
rect 44700 30690 44820 30810
rect 44940 30390 45060 30510
rect 46140 30690 46260 30810
rect 46620 27690 46740 27810
rect 45900 25590 46020 25710
rect 50940 32490 51060 32610
rect 47580 30090 47700 30210
rect 48780 27690 48900 27810
rect 48540 27390 48660 27510
rect 49020 27390 49140 27510
rect 46860 27090 46980 27210
rect 46860 26790 46980 26910
rect 46620 26490 46740 26610
rect 40140 25290 40260 25410
rect 41100 25290 41220 25410
rect 43740 25290 43860 25410
rect 46140 25290 46260 25410
rect 40380 24990 40500 25110
rect 40860 24990 40980 25110
rect 44460 24990 44580 25110
rect 40860 24390 40980 24510
rect 39660 24090 39780 24210
rect 39420 23790 39540 23910
rect 37020 22290 37140 22410
rect 36780 21390 36900 21510
rect 36780 21090 36900 21210
rect 38940 21690 39060 21810
rect 40620 23490 40740 23610
rect 39900 21690 40020 21810
rect 37500 20490 37620 20610
rect 37500 19890 37620 20010
rect 36540 19590 36660 19710
rect 37260 19590 37380 19710
rect 36540 19290 36660 19410
rect 36780 18390 36900 18510
rect 35820 16890 35940 17010
rect 39660 19290 39780 19410
rect 38940 18990 39060 19110
rect 39420 18990 39540 19110
rect 37260 17490 37380 17610
rect 35820 15690 35940 15810
rect 36300 15690 36420 15810
rect 34620 15390 34740 15510
rect 35340 15390 35460 15510
rect 32460 15090 32580 15210
rect 35100 15090 35220 15210
rect 36300 15390 36420 15510
rect 36060 15090 36180 15210
rect 37020 15090 37140 15210
rect 32700 14790 32820 14910
rect 33180 14790 33300 14910
rect 35580 14790 35700 14910
rect 36300 14790 36420 14910
rect 31980 13290 32100 13410
rect 31980 12990 32100 13110
rect 32460 12990 32580 13110
rect 32220 12390 32340 12510
rect 32220 12090 32340 12210
rect 32460 9090 32580 9210
rect 35820 14490 35940 14610
rect 34380 14190 34500 14310
rect 35340 13590 35460 13710
rect 32940 12990 33060 13110
rect 34620 13290 34740 13410
rect 34620 12990 34740 13110
rect 36060 12990 36180 13110
rect 34860 12690 34980 12810
rect 33180 9690 33300 9810
rect 36540 13290 36660 13410
rect 36780 12990 36900 13110
rect 36300 11790 36420 11910
rect 33660 9690 33780 9810
rect 32700 7590 32820 7710
rect 31740 6990 31860 7110
rect 32940 6990 33060 7110
rect 32220 6690 32340 6810
rect 24780 750 24900 870
rect 31500 6390 31620 6510
rect 35340 7590 35460 7710
rect 35100 7290 35220 7410
rect 33660 6690 33780 6810
rect 33180 6390 33300 6510
rect 34860 6390 34980 6510
rect 32460 6090 32580 6210
rect 38460 18390 38580 18510
rect 37980 15990 38100 16110
rect 37740 14790 37860 14910
rect 38220 15390 38340 15510
rect 40620 20790 40740 20910
rect 40380 19890 40500 20010
rect 42300 24090 42420 24210
rect 49980 27690 50100 27810
rect 48060 27090 48180 27210
rect 49020 26790 49140 26910
rect 47340 24990 47460 25110
rect 47820 23490 47940 23610
rect 42060 21690 42180 21810
rect 43980 21690 44100 21810
rect 42060 21390 42180 21510
rect 43740 21390 43860 21510
rect 42540 21090 42660 21210
rect 42300 20790 42420 20910
rect 42780 20790 42900 20910
rect 42300 19890 42420 20010
rect 43740 20790 43860 20910
rect 41580 19590 41700 19710
rect 42060 19590 42180 19710
rect 41100 19290 41220 19410
rect 41820 18990 41940 19110
rect 43500 18990 43620 19110
rect 45660 21090 45780 21210
rect 44940 20490 45060 20610
rect 45180 20190 45300 20310
rect 44700 18990 44820 19110
rect 43980 18690 44100 18810
rect 44460 18690 44580 18810
rect 40380 18390 40500 18510
rect 38940 18090 39060 18210
rect 40860 17790 40980 17910
rect 39420 15990 39540 16110
rect 38220 15090 38340 15210
rect 39420 14490 39540 14610
rect 43260 18390 43380 18510
rect 41340 15390 41460 15510
rect 42300 15690 42420 15810
rect 42300 15390 42420 15510
rect 41580 14790 41700 14910
rect 43020 15090 43140 15210
rect 42540 14190 42660 14310
rect 39420 12990 39540 13110
rect 40860 12990 40980 13110
rect 37980 12690 38100 12810
rect 37500 12390 37620 12510
rect 37260 9990 37380 10110
rect 36780 9690 36900 9810
rect 37500 9690 37620 9810
rect 38220 9690 38340 9810
rect 36540 7590 36660 7710
rect 36780 7290 36900 7410
rect 38700 12690 38820 12810
rect 38460 7590 38580 7710
rect 37260 7290 37380 7410
rect 39180 9390 39300 9510
rect 40620 12690 40740 12810
rect 41100 12390 41220 12510
rect 41580 12090 41700 12210
rect 41100 9990 41220 10110
rect 39420 9090 39540 9210
rect 39900 9390 40020 9510
rect 42060 9690 42180 9810
rect 40380 7590 40500 7710
rect 40860 7590 40980 7710
rect 38460 6990 38580 7110
rect 38940 6990 39060 7110
rect 38940 6690 39060 6810
rect 39420 6690 39540 6810
rect 37500 6390 37620 6510
rect 38460 6390 38580 6510
rect 36540 6090 36660 6210
rect 37020 6090 37140 6210
rect 43740 15690 43860 15810
rect 43260 14790 43380 14910
rect 44460 15690 44580 15810
rect 47340 21390 47460 21510
rect 49020 21990 49140 22110
rect 48060 21390 48180 21510
rect 46620 19890 46740 20010
rect 45420 18990 45540 19110
rect 47580 19890 47700 20010
rect 47580 19290 47700 19410
rect 48060 19290 48180 19410
rect 49980 20490 50100 20610
rect 46620 18690 46740 18810
rect 46620 18390 46740 18510
rect 49740 18390 49860 18510
rect 46860 17490 46980 17610
rect 46620 15690 46740 15810
rect 44700 15090 44820 15210
rect 45420 15090 45540 15210
rect 44460 12990 44580 13110
rect 45420 12990 45540 13110
rect 43260 12690 43380 12810
rect 43740 12690 43860 12810
rect 43740 11790 43860 11910
rect 42300 9090 42420 9210
rect 44460 12690 44580 12810
rect 44700 12390 44820 12510
rect 43980 9090 44100 9210
rect 42540 7890 42660 8010
rect 40860 6990 40980 7110
rect 46620 12690 46740 12810
rect 46620 12390 46740 12510
rect 44940 7590 45060 7710
rect 49260 15390 49380 15510
rect 49740 15390 49860 15510
rect 49500 15090 49620 15210
rect 48060 14790 48180 14910
rect 48300 13890 48420 14010
rect 47820 12390 47940 12510
rect 48300 12390 48420 12510
rect 48780 12390 48900 12510
rect 49260 12390 49380 12510
rect 46860 9690 46980 9810
rect 48540 12090 48660 12210
rect 47580 9090 47700 9210
rect 46620 7290 46740 7410
rect 44700 6990 44820 7110
rect 46620 6990 46740 7110
rect 48060 7890 48180 8010
rect 47340 7290 47460 7410
rect 44220 6690 44340 6810
rect 45420 6690 45540 6810
rect 46860 6690 46980 6810
rect 43980 6390 44100 6510
rect 47820 6390 47940 6510
rect 50220 12540 50340 12660
rect 50220 11490 50340 11610
rect 49500 9090 49620 9210
rect 50940 5190 51060 5310
rect 54540 11790 54660 11910
rect 54540 1020 54660 1140
<< metal3 >>
rect 18030 47025 18210 47040
rect 54480 47025 55350 47040
rect 18030 47010 55350 47025
rect 18030 46890 18060 47010
rect 18180 46890 55350 47010
rect 18030 46875 55350 46890
rect 18030 46860 18210 46875
rect 54480 46860 55350 46875
rect 15150 46725 15330 46740
rect 0 46710 15330 46725
rect 0 46590 15180 46710
rect 15300 46590 15330 46710
rect 0 46575 15330 46590
rect 15150 46560 15330 46575
rect 9390 44025 9570 44040
rect 22350 44025 22530 44040
rect 9390 44010 22530 44025
rect 9390 43890 9420 44010
rect 9540 43890 22380 44010
rect 22500 43890 22530 44010
rect 9390 43875 22530 43890
rect 9390 43860 9570 43875
rect 22350 43860 22530 43875
rect 7470 43725 7650 43740
rect 6285 43710 7650 43725
rect 6285 43590 7500 43710
rect 7620 43590 7650 43710
rect 6285 43575 7650 43590
rect 0 43425 6435 43575
rect 7470 43560 7650 43575
rect 18510 43725 18690 43740
rect 23310 43725 23490 43740
rect 18510 43710 23490 43725
rect 18510 43590 18540 43710
rect 18660 43590 23340 43710
rect 23460 43590 23490 43710
rect 18510 43575 23490 43590
rect 18510 43560 18690 43575
rect 23310 43560 23490 43575
rect 27630 43725 27810 43740
rect 28590 43725 28770 43740
rect 27630 43710 28770 43725
rect 27630 43590 27660 43710
rect 27780 43590 28620 43710
rect 28740 43590 28770 43710
rect 27630 43575 28770 43590
rect 27630 43560 27810 43575
rect 28590 43560 28770 43575
rect 36510 43725 36690 43740
rect 40110 43725 40290 43740
rect 36510 43710 40290 43725
rect 36510 43590 36540 43710
rect 36660 43590 40140 43710
rect 40260 43590 40290 43710
rect 36510 43575 40290 43590
rect 36510 43560 36690 43575
rect 40110 43560 40290 43575
rect 45630 43725 45810 43740
rect 46350 43725 46530 43740
rect 45630 43710 46530 43725
rect 45630 43590 45660 43710
rect 45780 43590 46380 43710
rect 46500 43590 46530 43710
rect 45630 43575 46530 43590
rect 45630 43560 45810 43575
rect 46350 43560 46530 43575
rect 12270 43425 12450 43440
rect 12990 43425 13170 43440
rect 12270 43410 13170 43425
rect 12270 43290 12300 43410
rect 12420 43290 13020 43410
rect 13140 43290 13170 43410
rect 12270 43275 13170 43290
rect 12270 43260 12450 43275
rect 12990 43260 13170 43275
rect 17070 43425 17250 43440
rect 18990 43425 19170 43440
rect 20190 43425 20370 43440
rect 17070 43410 20370 43425
rect 17070 43290 17100 43410
rect 17220 43290 19020 43410
rect 19140 43290 20220 43410
rect 20340 43290 20370 43410
rect 17070 43275 20370 43290
rect 17070 43260 17250 43275
rect 18990 43260 19170 43275
rect 20190 43260 20370 43275
rect 31470 43425 31650 43440
rect 40830 43425 41010 43440
rect 41310 43425 41490 43440
rect 42510 43425 42690 43440
rect 31470 43410 42690 43425
rect 31470 43290 31500 43410
rect 31620 43290 40860 43410
rect 40980 43290 41340 43410
rect 41460 43290 42540 43410
rect 42660 43290 42690 43410
rect 31470 43275 42690 43290
rect 31470 43260 31650 43275
rect 40830 43260 41010 43275
rect 41310 43260 41490 43275
rect 42510 43260 42690 43275
rect 6510 43125 6690 43140
rect 7230 43125 7410 43140
rect 6510 43110 7410 43125
rect 6510 42990 6540 43110
rect 6660 42990 7260 43110
rect 7380 42990 7410 43110
rect 6510 42975 7410 42990
rect 6510 42960 6690 42975
rect 7230 42960 7410 42975
rect 8670 43125 8850 43140
rect 10350 43125 10530 43140
rect 8670 43110 10530 43125
rect 8670 42990 8700 43110
rect 8820 42990 10380 43110
rect 10500 42990 10530 43110
rect 8670 42975 10530 42990
rect 8670 42960 8850 42975
rect 10350 42960 10530 42975
rect 10830 43125 11010 43140
rect 11310 43125 11490 43140
rect 10830 43110 11490 43125
rect 10830 42990 10860 43110
rect 10980 42990 11340 43110
rect 11460 42990 11490 43110
rect 10830 42975 11490 42990
rect 10830 42960 11010 42975
rect 11310 42960 11490 42975
rect 13710 43125 13890 43140
rect 14670 43125 14850 43140
rect 13710 43110 14850 43125
rect 13710 42990 13740 43110
rect 13860 42990 14700 43110
rect 14820 42990 14850 43110
rect 13710 42975 14850 42990
rect 13710 42960 13890 42975
rect 14670 42960 14850 42975
rect 28110 43125 28290 43140
rect 28830 43125 29010 43140
rect 32190 43125 32370 43140
rect 28110 43110 32370 43125
rect 28110 42990 28140 43110
rect 28260 42990 28860 43110
rect 28980 42990 32220 43110
rect 32340 42990 32370 43110
rect 28110 42975 32370 42990
rect 28110 42960 28290 42975
rect 28830 42960 29010 42975
rect 32190 42960 32370 42975
rect 34590 43125 34770 43140
rect 35070 43125 35250 43140
rect 34590 43110 35250 43125
rect 34590 42990 34620 43110
rect 34740 42990 35100 43110
rect 35220 42990 35250 43110
rect 34590 42975 35250 42990
rect 34590 42960 34770 42975
rect 35070 42960 35250 42975
rect 37230 43125 37410 43140
rect 38430 43125 38610 43140
rect 37230 43110 38610 43125
rect 37230 42990 37260 43110
rect 37380 42990 38460 43110
rect 38580 42990 38610 43110
rect 37230 42975 38610 42990
rect 37230 42960 37410 42975
rect 38430 42960 38610 42975
rect 44190 43125 44370 43140
rect 44670 43125 44850 43140
rect 45390 43125 45570 43140
rect 44190 43110 45570 43125
rect 44190 42990 44220 43110
rect 44340 42990 44700 43110
rect 44820 42990 45420 43110
rect 45540 42990 45570 43110
rect 44190 42975 45570 42990
rect 44190 42960 44370 42975
rect 44670 42960 44850 42975
rect 45390 42960 45570 42975
rect 6750 42825 6930 42840
rect 9630 42825 9810 42840
rect 6750 42810 9810 42825
rect 6750 42690 6780 42810
rect 6900 42690 9660 42810
rect 9780 42690 9810 42810
rect 6750 42675 9810 42690
rect 6750 42660 6930 42675
rect 9630 42660 9810 42675
rect 13950 42825 14130 42840
rect 15870 42825 16050 42840
rect 13950 42810 16050 42825
rect 13950 42690 13980 42810
rect 14100 42690 15900 42810
rect 16020 42690 16050 42810
rect 13950 42675 16050 42690
rect 13950 42660 14130 42675
rect 15870 42660 16050 42675
rect 17310 42825 17490 42840
rect 20670 42825 20850 42840
rect 17310 42810 20850 42825
rect 17310 42690 17340 42810
rect 17460 42690 20700 42810
rect 20820 42690 20850 42810
rect 17310 42675 20850 42690
rect 17310 42660 17490 42675
rect 20670 42660 20850 42675
rect 30510 42825 30690 42840
rect 31230 42825 31410 42840
rect 30510 42810 31410 42825
rect 30510 42690 30540 42810
rect 30660 42690 31260 42810
rect 31380 42690 31410 42810
rect 30510 42675 31410 42690
rect 30510 42660 30690 42675
rect 31230 42660 31410 42675
rect 31950 42825 32130 42840
rect 32430 42825 32610 42840
rect 33630 42825 33810 42840
rect 36510 42825 36690 42840
rect 31950 42810 36690 42825
rect 31950 42690 31980 42810
rect 32100 42690 32460 42810
rect 32580 42690 33660 42810
rect 33780 42690 36540 42810
rect 36660 42690 36690 42810
rect 31950 42675 36690 42690
rect 31950 42660 32130 42675
rect 32430 42660 32610 42675
rect 33630 42660 33810 42675
rect 36510 42660 36690 42675
rect 44430 42825 44610 42840
rect 44910 42825 45090 42840
rect 44430 42810 45090 42825
rect 44430 42690 44460 42810
rect 44580 42690 44940 42810
rect 45060 42690 45090 42810
rect 44430 42675 45090 42690
rect 44430 42660 44610 42675
rect 44910 42660 45090 42675
rect 5550 42525 5730 42540
rect 6510 42525 6690 42540
rect 5550 42510 6690 42525
rect 5550 42390 5580 42510
rect 5700 42390 6540 42510
rect 6660 42390 6690 42510
rect 5550 42375 6690 42390
rect 5550 42360 5730 42375
rect 6510 42360 6690 42375
rect 7710 42525 7890 42540
rect 8430 42525 8610 42540
rect 7710 42510 8610 42525
rect 7710 42390 7740 42510
rect 7860 42390 8460 42510
rect 8580 42390 8610 42510
rect 7710 42375 8610 42390
rect 7710 42360 7890 42375
rect 8430 42360 8610 42375
rect 8910 42525 9090 42540
rect 9630 42525 9810 42540
rect 8910 42510 9810 42525
rect 8910 42390 8940 42510
rect 9060 42390 9660 42510
rect 9780 42390 9810 42510
rect 8910 42375 9810 42390
rect 8910 42360 9090 42375
rect 9630 42360 9810 42375
rect 15870 42525 16050 42540
rect 18030 42525 18210 42540
rect 15870 42510 18210 42525
rect 15870 42390 15900 42510
rect 16020 42390 18060 42510
rect 18180 42390 18210 42510
rect 15870 42375 18210 42390
rect 15870 42360 16050 42375
rect 18030 42360 18210 42375
rect 19230 42525 19410 42540
rect 19710 42525 19890 42540
rect 19230 42510 19890 42525
rect 19230 42390 19260 42510
rect 19380 42390 19740 42510
rect 19860 42390 19890 42510
rect 19230 42375 19890 42390
rect 19230 42360 19410 42375
rect 19710 42360 19890 42375
rect 24990 42525 25170 42540
rect 25950 42525 26130 42540
rect 24990 42510 26130 42525
rect 24990 42390 25020 42510
rect 25140 42390 25980 42510
rect 26100 42390 26130 42510
rect 24990 42375 26130 42390
rect 24990 42360 25170 42375
rect 25950 42360 26130 42375
rect 27870 42525 28050 42540
rect 29550 42525 29730 42540
rect 27870 42510 29730 42525
rect 27870 42390 27900 42510
rect 28020 42390 29580 42510
rect 29700 42390 29730 42510
rect 27870 42375 29730 42390
rect 27870 42360 28050 42375
rect 29550 42360 29730 42375
rect 31470 42525 31650 42540
rect 32190 42525 32370 42540
rect 31470 42510 32370 42525
rect 31470 42390 31500 42510
rect 31620 42390 32220 42510
rect 32340 42390 32370 42510
rect 31470 42375 32370 42390
rect 31470 42360 31650 42375
rect 32190 42360 32370 42375
rect 46110 42525 46290 42540
rect 47310 42525 47490 42540
rect 46110 42510 47490 42525
rect 46110 42390 46140 42510
rect 46260 42390 47340 42510
rect 47460 42390 47490 42510
rect 46110 42375 47490 42390
rect 46110 42360 46290 42375
rect 47310 42360 47490 42375
rect 25710 42225 25890 42240
rect 27150 42225 27330 42240
rect 25710 42210 27330 42225
rect 25710 42090 25740 42210
rect 25860 42090 27180 42210
rect 27300 42090 27330 42210
rect 25710 42075 27330 42090
rect 25710 42060 25890 42075
rect 27150 42060 27330 42075
rect 31230 42225 31410 42240
rect 33150 42225 33330 42240
rect 31230 42210 33330 42225
rect 31230 42090 31260 42210
rect 31380 42090 33180 42210
rect 33300 42090 33330 42210
rect 31230 42075 33330 42090
rect 31230 42060 31410 42075
rect 33150 42060 33330 42075
rect 44910 42225 45090 42240
rect 46590 42225 46770 42240
rect 44910 42210 46770 42225
rect 44910 42090 44940 42210
rect 45060 42090 46620 42210
rect 46740 42090 46770 42210
rect 44910 42075 46770 42090
rect 44910 42060 45090 42075
rect 46590 42060 46770 42075
rect 43470 41925 43650 41940
rect 48750 41925 48930 41940
rect 43470 41910 48930 41925
rect 43470 41790 43500 41910
rect 43620 41790 48780 41910
rect 48900 41790 48930 41910
rect 43470 41775 48930 41790
rect 43470 41760 43650 41775
rect 48750 41760 48930 41775
rect 45630 41625 45810 41640
rect 46830 41625 47010 41640
rect 45630 41610 47010 41625
rect 45630 41490 45660 41610
rect 45780 41490 46860 41610
rect 46980 41490 47010 41610
rect 45630 41475 47010 41490
rect 45630 41460 45810 41475
rect 46830 41460 47010 41475
rect 15630 41325 15810 41340
rect 28830 41325 29010 41340
rect 15630 41310 29010 41325
rect 15630 41190 15660 41310
rect 15780 41190 28860 41310
rect 28980 41190 29010 41310
rect 15630 41175 29010 41190
rect 15630 41160 15810 41175
rect 28830 41160 29010 41175
rect 22590 41025 22770 41040
rect 24030 41025 24210 41040
rect 22590 41010 24210 41025
rect 22590 40890 22620 41010
rect 22740 40890 24060 41010
rect 24180 40890 24210 41010
rect 22590 40875 24210 40890
rect 22590 40860 22770 40875
rect 24030 40860 24210 40875
rect 26190 40725 26370 40740
rect 34110 40725 34290 40740
rect 26190 40710 34290 40725
rect 26190 40590 26220 40710
rect 26340 40590 34140 40710
rect 34260 40590 34290 40710
rect 26190 40575 34290 40590
rect 26190 40560 26370 40575
rect 34110 40560 34290 40575
rect 11310 40125 11490 40140
rect 12750 40125 12930 40140
rect 14430 40125 14610 40140
rect 11310 40110 14610 40125
rect 11310 39990 11340 40110
rect 11460 39990 12780 40110
rect 12900 39990 14460 40110
rect 14580 39990 14610 40110
rect 11310 39975 14610 39990
rect 11310 39960 11490 39975
rect 12750 39960 12930 39975
rect 14430 39960 14610 39975
rect 46830 39825 47010 39840
rect 49230 39825 49410 39840
rect 46830 39810 49410 39825
rect 46830 39690 46860 39810
rect 46980 39690 49260 39810
rect 49380 39690 49410 39810
rect 46830 39675 49410 39690
rect 46830 39660 47010 39675
rect 49230 39660 49410 39675
rect 9630 39525 9810 39540
rect 12990 39525 13170 39540
rect 9630 39510 13170 39525
rect 9630 39390 9660 39510
rect 9780 39390 13020 39510
rect 13140 39390 13170 39510
rect 9630 39375 13170 39390
rect 9630 39360 9810 39375
rect 12990 39360 13170 39375
rect 19470 39525 19650 39540
rect 21390 39525 21570 39540
rect 19470 39510 21570 39525
rect 19470 39390 19500 39510
rect 19620 39390 21420 39510
rect 21540 39390 21570 39510
rect 19470 39375 21570 39390
rect 19470 39360 19650 39375
rect 21390 39360 21570 39375
rect 24030 39525 24210 39540
rect 27150 39525 27330 39540
rect 24030 39510 27330 39525
rect 24030 39390 24060 39510
rect 24180 39390 27180 39510
rect 27300 39390 27330 39510
rect 24030 39375 27330 39390
rect 24030 39360 24210 39375
rect 27150 39360 27330 39375
rect 39150 39525 39330 39540
rect 40830 39525 41010 39540
rect 41550 39525 41730 39540
rect 42270 39525 42450 39540
rect 39150 39510 42450 39525
rect 39150 39390 39180 39510
rect 39300 39390 40860 39510
rect 40980 39390 41580 39510
rect 41700 39390 42300 39510
rect 42420 39390 42450 39510
rect 39150 39375 42450 39390
rect 39150 39360 39330 39375
rect 40830 39360 41010 39375
rect 41550 39360 41730 39375
rect 42270 39360 42450 39375
rect 45870 39525 46050 39540
rect 46350 39525 46530 39540
rect 45870 39510 46530 39525
rect 45870 39390 45900 39510
rect 46020 39390 46380 39510
rect 46500 39390 46530 39510
rect 45870 39375 46530 39390
rect 45870 39360 46050 39375
rect 46350 39360 46530 39375
rect 6030 39225 6210 39240
rect 7470 39225 7650 39240
rect 6030 39210 7650 39225
rect 6030 39090 6060 39210
rect 6180 39090 7500 39210
rect 7620 39090 7650 39210
rect 6030 39075 7650 39090
rect 6030 39060 6210 39075
rect 7470 39060 7650 39075
rect 13230 39225 13410 39240
rect 14190 39225 14370 39240
rect 13230 39210 14370 39225
rect 13230 39090 13260 39210
rect 13380 39090 14220 39210
rect 14340 39090 14370 39210
rect 13230 39075 14370 39090
rect 13230 39060 13410 39075
rect 14190 39060 14370 39075
rect 18270 39225 18450 39240
rect 18750 39225 18930 39240
rect 20910 39225 21090 39240
rect 18270 39210 21090 39225
rect 18270 39090 18300 39210
rect 18420 39090 18780 39210
rect 18900 39090 20940 39210
rect 21060 39090 21090 39210
rect 18270 39075 21090 39090
rect 18270 39060 18450 39075
rect 18750 39060 18930 39075
rect 20910 39060 21090 39075
rect 23790 39225 23970 39240
rect 24270 39225 24450 39240
rect 27150 39225 27330 39240
rect 23790 39210 27330 39225
rect 23790 39090 23820 39210
rect 23940 39090 24300 39210
rect 24420 39090 27180 39210
rect 27300 39090 27330 39210
rect 23790 39075 27330 39090
rect 23790 39060 23970 39075
rect 24270 39060 24450 39075
rect 27150 39060 27330 39075
rect 33390 39225 33570 39240
rect 35070 39225 35250 39240
rect 35550 39225 35730 39240
rect 36030 39225 36210 39240
rect 33390 39210 36210 39225
rect 33390 39090 33420 39210
rect 33540 39090 35100 39210
rect 35220 39090 35580 39210
rect 35700 39090 36060 39210
rect 36180 39090 36210 39210
rect 33390 39075 36210 39090
rect 33390 39060 33570 39075
rect 35070 39060 35250 39075
rect 35550 39060 35730 39075
rect 36030 39060 36210 39075
rect 38910 39225 39090 39240
rect 39870 39225 40050 39240
rect 43710 39225 43890 39240
rect 45150 39225 45330 39240
rect 38910 39210 45330 39225
rect 38910 39090 38940 39210
rect 39060 39090 39900 39210
rect 40020 39090 43740 39210
rect 43860 39090 45180 39210
rect 45300 39090 45330 39210
rect 38910 39075 45330 39090
rect 38910 39060 39090 39075
rect 39870 39060 40050 39075
rect 43710 39060 43890 39075
rect 45150 39060 45330 39075
rect 47070 39225 47250 39240
rect 48030 39225 48210 39240
rect 47070 39210 48210 39225
rect 47070 39090 47100 39210
rect 47220 39090 48060 39210
rect 48180 39090 48210 39210
rect 47070 39075 48210 39090
rect 47070 39060 47250 39075
rect 48030 39060 48210 39075
rect 2430 38925 2610 38940
rect 17550 38925 17730 38940
rect 2430 38910 17730 38925
rect 2430 38790 2460 38910
rect 2580 38790 17580 38910
rect 17700 38790 17730 38910
rect 2430 38775 17730 38790
rect 2430 38760 2610 38775
rect 17550 38760 17730 38775
rect 21870 38925 22050 38940
rect 23550 38925 23730 38940
rect 24750 38925 24930 38940
rect 21870 38910 24930 38925
rect 21870 38790 21900 38910
rect 22020 38790 23580 38910
rect 23700 38790 24780 38910
rect 24900 38790 24930 38910
rect 21870 38775 24930 38790
rect 21870 38760 22050 38775
rect 23550 38760 23730 38775
rect 24750 38760 24930 38775
rect 25710 38925 25890 38940
rect 28110 38925 28290 38940
rect 33390 38925 33570 38940
rect 25710 38910 33570 38925
rect 25710 38790 25740 38910
rect 25860 38790 28140 38910
rect 28260 38790 33420 38910
rect 33540 38790 33570 38910
rect 25710 38775 33570 38790
rect 25710 38760 25890 38775
rect 28110 38760 28290 38775
rect 33390 38760 33570 38775
rect 38190 38925 38370 38940
rect 40830 38925 41010 38940
rect 38190 38910 41010 38925
rect 38190 38790 38220 38910
rect 38340 38790 40860 38910
rect 40980 38790 41010 38910
rect 38190 38775 41010 38790
rect 38190 38760 38370 38775
rect 40830 38760 41010 38775
rect 47790 38925 47970 38940
rect 49710 38925 49890 38940
rect 47790 38910 49890 38925
rect 47790 38790 47820 38910
rect 47940 38790 49740 38910
rect 49860 38790 49890 38910
rect 47790 38775 49890 38790
rect 47790 38760 47970 38775
rect 49710 38760 49890 38775
rect 16110 38625 16290 38640
rect 30750 38625 30930 38640
rect 16110 38610 30930 38625
rect 16110 38490 16140 38610
rect 16260 38490 30780 38610
rect 30900 38490 30930 38610
rect 16110 38475 30930 38490
rect 16110 38460 16290 38475
rect 30750 38460 30930 38475
rect 37470 38625 37650 38640
rect 40590 38625 40770 38640
rect 37470 38610 40770 38625
rect 37470 38490 37500 38610
rect 37620 38490 40620 38610
rect 40740 38490 40770 38610
rect 37470 38475 40770 38490
rect 37470 38460 37650 38475
rect 40590 38460 40770 38475
rect 43710 38625 43890 38640
rect 45390 38625 45570 38640
rect 43710 38610 45570 38625
rect 43710 38490 43740 38610
rect 43860 38490 45420 38610
rect 45540 38490 45570 38610
rect 43710 38475 45570 38490
rect 43710 38460 43890 38475
rect 45390 38460 45570 38475
rect 5310 38175 5490 38190
rect 0 38160 5490 38175
rect 0 38040 5340 38160
rect 5460 38040 5490 38160
rect 0 38025 5490 38040
rect 5310 38010 5490 38025
rect 2670 37725 2850 37740
rect 12270 37725 12450 37740
rect 2670 37710 12450 37725
rect 2670 37590 2700 37710
rect 2820 37590 12300 37710
rect 12420 37590 12450 37710
rect 2670 37575 12450 37590
rect 2670 37560 2850 37575
rect 12270 37560 12450 37575
rect 31230 37725 31410 37740
rect 32910 37725 33090 37740
rect 31230 37710 33090 37725
rect 31230 37590 31260 37710
rect 31380 37590 32940 37710
rect 33060 37590 33090 37710
rect 31230 37575 33090 37590
rect 31230 37560 31410 37575
rect 32910 37560 33090 37575
rect 35790 37725 35970 37740
rect 39390 37725 39570 37740
rect 35790 37710 39570 37725
rect 35790 37590 35820 37710
rect 35940 37590 39420 37710
rect 39540 37590 39570 37710
rect 35790 37575 39570 37590
rect 35790 37560 35970 37575
rect 39390 37560 39570 37575
rect 2670 37425 2850 37440
rect 10830 37425 11010 37440
rect 2670 37410 11010 37425
rect 2670 37290 2700 37410
rect 2820 37290 10860 37410
rect 10980 37290 11010 37410
rect 2670 37275 11010 37290
rect 2670 37260 2850 37275
rect 10830 37260 11010 37275
rect 12030 37425 12210 37440
rect 17070 37425 17250 37440
rect 12030 37410 17250 37425
rect 12030 37290 12060 37410
rect 12180 37290 17100 37410
rect 17220 37290 17250 37410
rect 12030 37275 17250 37290
rect 12030 37260 12210 37275
rect 17070 37260 17250 37275
rect 22350 37425 22530 37440
rect 24270 37425 24450 37440
rect 22350 37410 24450 37425
rect 22350 37290 22380 37410
rect 22500 37290 24300 37410
rect 24420 37290 24450 37410
rect 22350 37275 24450 37290
rect 22350 37260 22530 37275
rect 24270 37260 24450 37275
rect 30030 37425 30210 37440
rect 30990 37425 31170 37440
rect 30030 37410 31170 37425
rect 30030 37290 30060 37410
rect 30180 37290 31020 37410
rect 31140 37290 31170 37410
rect 30030 37275 31170 37290
rect 30030 37260 30210 37275
rect 30990 37260 31170 37275
rect 32670 37425 32850 37440
rect 36990 37425 37170 37440
rect 32670 37410 37170 37425
rect 32670 37290 32700 37410
rect 32820 37290 37020 37410
rect 37140 37290 37170 37410
rect 32670 37275 37170 37290
rect 32670 37260 32850 37275
rect 36990 37260 37170 37275
rect 40350 37425 40530 37440
rect 43950 37425 44130 37440
rect 46590 37425 46770 37440
rect 40350 37410 46770 37425
rect 40350 37290 40380 37410
rect 40500 37290 43980 37410
rect 44100 37290 46620 37410
rect 46740 37290 46770 37410
rect 40350 37275 46770 37290
rect 40350 37260 40530 37275
rect 43950 37260 44130 37275
rect 46590 37260 46770 37275
rect 6750 37125 6930 37140
rect 7230 37125 7410 37140
rect 6750 37110 7410 37125
rect 6750 36990 6780 37110
rect 6900 36990 7260 37110
rect 7380 36990 7410 37110
rect 6750 36975 7410 36990
rect 6750 36960 6930 36975
rect 7230 36960 7410 36975
rect 10830 37125 11010 37140
rect 12990 37125 13170 37140
rect 10830 37110 13170 37125
rect 10830 36990 10860 37110
rect 10980 36990 13020 37110
rect 13140 36990 13170 37110
rect 10830 36975 13170 36990
rect 10830 36960 11010 36975
rect 12990 36960 13170 36975
rect 14670 37125 14850 37140
rect 15390 37125 15570 37140
rect 16350 37125 16530 37140
rect 18510 37125 18690 37140
rect 14670 37110 18690 37125
rect 14670 36990 14700 37110
rect 14820 36990 15420 37110
rect 15540 36990 16380 37110
rect 16500 36990 18540 37110
rect 18660 36990 18690 37110
rect 14670 36975 18690 36990
rect 14670 36960 14850 36975
rect 15390 36960 15570 36975
rect 16350 36960 16530 36975
rect 18510 36960 18690 36975
rect 20910 37125 21090 37140
rect 21390 37125 21570 37140
rect 20910 37110 21570 37125
rect 20910 36990 20940 37110
rect 21060 36990 21420 37110
rect 21540 36990 21570 37110
rect 20910 36975 21570 36990
rect 20910 36960 21090 36975
rect 21390 36960 21570 36975
rect 23790 37125 23970 37140
rect 24990 37125 25170 37140
rect 25710 37125 25890 37140
rect 27870 37125 28050 37140
rect 28350 37125 28530 37140
rect 23790 37110 25890 37125
rect 23790 36990 23820 37110
rect 23940 36990 25020 37110
rect 25140 36990 25740 37110
rect 25860 36990 25890 37110
rect 23790 36975 25890 36990
rect 23790 36960 23970 36975
rect 24990 36960 25170 36975
rect 25710 36960 25890 36975
rect 27405 37110 28530 37125
rect 27405 36990 27900 37110
rect 28020 36990 28380 37110
rect 28500 36990 28530 37110
rect 27405 36975 28530 36990
rect 10830 36825 11010 36840
rect 11310 36825 11490 36840
rect 10830 36810 11490 36825
rect 10830 36690 10860 36810
rect 10980 36690 11340 36810
rect 11460 36690 11490 36810
rect 10830 36675 11490 36690
rect 10830 36660 11010 36675
rect 11310 36660 11490 36675
rect 19470 36825 19650 36840
rect 27405 36825 27555 36975
rect 27870 36960 28050 36975
rect 28350 36960 28530 36975
rect 32910 37125 33090 37140
rect 35070 37125 35250 37140
rect 32910 37110 35250 37125
rect 32910 36990 32940 37110
rect 33060 36990 35100 37110
rect 35220 36990 35250 37110
rect 32910 36975 35250 36990
rect 32910 36960 33090 36975
rect 35070 36960 35250 36975
rect 43230 37125 43410 37140
rect 43710 37125 43890 37140
rect 43230 37110 43890 37125
rect 43230 36990 43260 37110
rect 43380 36990 43740 37110
rect 43860 36990 43890 37110
rect 43230 36975 43890 36990
rect 43230 36960 43410 36975
rect 43710 36960 43890 36975
rect 44670 37125 44850 37140
rect 45390 37125 45570 37140
rect 48030 37125 48210 37140
rect 44670 37110 48210 37125
rect 44670 36990 44700 37110
rect 44820 36990 45420 37110
rect 45540 36990 48060 37110
rect 48180 36990 48210 37110
rect 44670 36975 48210 36990
rect 44670 36960 44850 36975
rect 45390 36960 45570 36975
rect 48030 36960 48210 36975
rect 19470 36810 27555 36825
rect 19470 36690 19500 36810
rect 19620 36690 27555 36810
rect 19470 36675 27555 36690
rect 31950 36825 32130 36840
rect 32430 36825 32610 36840
rect 31950 36810 32610 36825
rect 31950 36690 31980 36810
rect 32100 36690 32460 36810
rect 32580 36690 32610 36810
rect 31950 36675 32610 36690
rect 19470 36660 19650 36675
rect 31950 36660 32130 36675
rect 32430 36660 32610 36675
rect 42270 36825 42450 36840
rect 42750 36825 42930 36840
rect 42270 36810 42930 36825
rect 42270 36690 42300 36810
rect 42420 36690 42780 36810
rect 42900 36690 42930 36810
rect 42270 36675 42930 36690
rect 42270 36660 42450 36675
rect 42750 36660 42930 36675
rect 47790 36825 47970 36840
rect 49710 36825 49890 36840
rect 47790 36810 49890 36825
rect 47790 36690 47820 36810
rect 47940 36690 49740 36810
rect 49860 36690 49890 36810
rect 47790 36675 49890 36690
rect 47790 36660 47970 36675
rect 49710 36660 49890 36675
rect 50430 36675 50610 36690
rect 55200 36675 55350 36690
rect 50430 36660 55350 36675
rect 50430 36540 50460 36660
rect 50580 36540 55350 36660
rect 5550 36525 5730 36540
rect 6990 36525 7170 36540
rect 5550 36510 7170 36525
rect 5550 36390 5580 36510
rect 5700 36390 7020 36510
rect 7140 36390 7170 36510
rect 5550 36375 7170 36390
rect 5550 36360 5730 36375
rect 6990 36360 7170 36375
rect 8190 36525 8370 36540
rect 9150 36525 9330 36540
rect 8190 36510 9330 36525
rect 8190 36390 8220 36510
rect 8340 36390 9180 36510
rect 9300 36390 9330 36510
rect 8190 36375 9330 36390
rect 8190 36360 8370 36375
rect 9150 36360 9330 36375
rect 14910 36525 15090 36540
rect 16110 36525 16290 36540
rect 14910 36510 16290 36525
rect 14910 36390 14940 36510
rect 15060 36390 16140 36510
rect 16260 36390 16290 36510
rect 14910 36375 16290 36390
rect 14910 36360 15090 36375
rect 16110 36360 16290 36375
rect 19950 36525 20130 36540
rect 21390 36525 21570 36540
rect 19950 36510 21570 36525
rect 19950 36390 19980 36510
rect 20100 36390 21420 36510
rect 21540 36390 21570 36510
rect 19950 36375 21570 36390
rect 19950 36360 20130 36375
rect 21390 36360 21570 36375
rect 26190 36525 26370 36540
rect 27150 36525 27330 36540
rect 26190 36510 27330 36525
rect 26190 36390 26220 36510
rect 26340 36390 27180 36510
rect 27300 36390 27330 36510
rect 26190 36375 27330 36390
rect 26190 36360 26370 36375
rect 27150 36360 27330 36375
rect 31230 36525 31410 36540
rect 31710 36525 31890 36540
rect 31230 36510 31890 36525
rect 31230 36390 31260 36510
rect 31380 36390 31740 36510
rect 31860 36390 31890 36510
rect 31230 36375 31890 36390
rect 31230 36360 31410 36375
rect 31710 36360 31890 36375
rect 33150 36525 33330 36540
rect 33630 36525 33810 36540
rect 33150 36510 33810 36525
rect 33150 36390 33180 36510
rect 33300 36390 33660 36510
rect 33780 36390 33810 36510
rect 33150 36375 33810 36390
rect 33150 36360 33330 36375
rect 33630 36360 33810 36375
rect 34350 36525 34530 36540
rect 39390 36525 39570 36540
rect 34350 36510 39570 36525
rect 34350 36390 34380 36510
rect 34500 36390 39420 36510
rect 39540 36390 39570 36510
rect 34350 36375 39570 36390
rect 34350 36360 34530 36375
rect 39390 36360 39570 36375
rect 47550 36525 47730 36540
rect 48270 36525 48450 36540
rect 49230 36525 49410 36540
rect 47550 36510 49410 36525
rect 50430 36525 55350 36540
rect 50430 36510 50610 36525
rect 55200 36510 55350 36525
rect 47550 36390 47580 36510
rect 47700 36390 48300 36510
rect 48420 36390 49260 36510
rect 49380 36390 49410 36510
rect 47550 36375 49410 36390
rect 47550 36360 47730 36375
rect 48270 36360 48450 36375
rect 49230 36360 49410 36375
rect 10110 36225 10290 36240
rect 16110 36225 16290 36240
rect 10110 36210 16290 36225
rect 10110 36090 10140 36210
rect 10260 36090 16140 36210
rect 16260 36090 16290 36210
rect 10110 36075 16290 36090
rect 10110 36060 10290 36075
rect 16110 36060 16290 36075
rect 21390 36225 21570 36240
rect 23070 36225 23250 36240
rect 28350 36225 28530 36240
rect 21390 36210 28530 36225
rect 21390 36090 21420 36210
rect 21540 36090 23100 36210
rect 23220 36090 28380 36210
rect 28500 36090 28530 36210
rect 21390 36075 28530 36090
rect 21390 36060 21570 36075
rect 23070 36060 23250 36075
rect 28350 36060 28530 36075
rect 28830 36225 29010 36240
rect 35070 36225 35250 36240
rect 28830 36210 35250 36225
rect 28830 36090 28860 36210
rect 28980 36090 35100 36210
rect 35220 36090 35250 36210
rect 28830 36075 35250 36090
rect 28830 36060 29010 36075
rect 35070 36060 35250 36075
rect 36270 36225 36450 36240
rect 41310 36225 41490 36240
rect 42270 36225 42450 36240
rect 36270 36210 42450 36225
rect 36270 36090 36300 36210
rect 36420 36090 41340 36210
rect 41460 36090 42300 36210
rect 42420 36090 42450 36210
rect 36270 36075 42450 36090
rect 36270 36060 36450 36075
rect 41310 36060 41490 36075
rect 42270 36060 42450 36075
rect 22830 35925 23010 35940
rect 29550 35925 29730 35940
rect 35310 35925 35490 35940
rect 22830 35910 35490 35925
rect 22830 35790 22860 35910
rect 22980 35790 29580 35910
rect 29700 35790 35340 35910
rect 35460 35790 35490 35910
rect 22830 35775 35490 35790
rect 22830 35760 23010 35775
rect 29550 35760 29730 35775
rect 35310 35760 35490 35775
rect 40350 35625 40530 35640
rect 43230 35625 43410 35640
rect 40350 35610 43410 35625
rect 40350 35490 40380 35610
rect 40500 35490 43260 35610
rect 43380 35490 43410 35610
rect 40350 35475 43410 35490
rect 40350 35460 40530 35475
rect 43230 35460 43410 35475
rect 28350 35325 28530 35340
rect 50430 35325 50610 35340
rect 28350 35310 50610 35325
rect 28350 35190 28380 35310
rect 28500 35190 50460 35310
rect 50580 35190 50610 35310
rect 28350 35175 50610 35190
rect 28350 35160 28530 35175
rect 50430 35160 50610 35175
rect 36270 35025 36450 35040
rect 46830 35025 47010 35040
rect 36270 35010 47010 35025
rect 36270 34890 36300 35010
rect 36420 34890 46860 35010
rect 46980 34890 47010 35010
rect 36270 34875 47010 34890
rect 36270 34860 36450 34875
rect 46830 34860 47010 34875
rect 34830 34725 35010 34740
rect 37230 34725 37410 34740
rect 34830 34710 37410 34725
rect 34830 34590 34860 34710
rect 34980 34590 37260 34710
rect 37380 34590 37410 34710
rect 34830 34575 37410 34590
rect 34830 34560 35010 34575
rect 37230 34560 37410 34575
rect 15150 34425 15330 34440
rect 18750 34425 18930 34440
rect 15150 34410 18930 34425
rect 15150 34290 15180 34410
rect 15300 34290 18780 34410
rect 18900 34290 18930 34410
rect 15150 34275 18930 34290
rect 15150 34260 15330 34275
rect 18750 34260 18930 34275
rect 24750 34425 24930 34440
rect 33390 34425 33570 34440
rect 24750 34410 33570 34425
rect 24750 34290 24780 34410
rect 24900 34290 33420 34410
rect 33540 34290 33570 34410
rect 24750 34275 33570 34290
rect 24750 34260 24930 34275
rect 33390 34260 33570 34275
rect 12750 34125 12930 34140
rect 19710 34125 19890 34140
rect 12750 34110 19890 34125
rect 12750 33990 12780 34110
rect 12900 33990 19740 34110
rect 19860 33990 19890 34110
rect 12750 33975 19890 33990
rect 12750 33960 12930 33975
rect 19710 33960 19890 33975
rect 30510 34125 30690 34140
rect 32670 34125 32850 34140
rect 30510 34110 32850 34125
rect 30510 33990 30540 34110
rect 30660 33990 32700 34110
rect 32820 33990 32850 34110
rect 30510 33975 32850 33990
rect 30510 33960 30690 33975
rect 32670 33960 32850 33975
rect 35070 34125 35250 34140
rect 36270 34125 36450 34140
rect 35070 34110 36450 34125
rect 35070 33990 35100 34110
rect 35220 33990 36300 34110
rect 36420 33990 36450 34110
rect 35070 33975 36450 33990
rect 35070 33960 35250 33975
rect 36270 33960 36450 33975
rect 41550 34125 41730 34140
rect 42030 34125 42210 34140
rect 41550 34110 42210 34125
rect 41550 33990 41580 34110
rect 41700 33990 42060 34110
rect 42180 33990 42210 34110
rect 41550 33975 42210 33990
rect 41550 33960 41730 33975
rect 42030 33960 42210 33975
rect 7230 33825 7410 33840
rect 7710 33825 7890 33840
rect 7230 33810 7890 33825
rect 7230 33690 7260 33810
rect 7380 33690 7740 33810
rect 7860 33690 7890 33810
rect 7230 33675 7890 33690
rect 7230 33660 7410 33675
rect 7710 33660 7890 33675
rect 17310 33825 17490 33840
rect 18510 33825 18690 33840
rect 21150 33825 21330 33840
rect 17310 33810 21330 33825
rect 17310 33690 17340 33810
rect 17460 33690 18540 33810
rect 18660 33690 21180 33810
rect 21300 33690 21330 33810
rect 17310 33675 21330 33690
rect 17310 33660 17490 33675
rect 18510 33660 18690 33675
rect 21150 33660 21330 33675
rect 24510 33825 24690 33840
rect 25230 33825 25410 33840
rect 24510 33810 25410 33825
rect 24510 33690 24540 33810
rect 24660 33690 25260 33810
rect 25380 33690 25410 33810
rect 24510 33675 25410 33690
rect 24510 33660 24690 33675
rect 25230 33660 25410 33675
rect 31710 33825 31890 33840
rect 32670 33825 32850 33840
rect 31710 33810 32850 33825
rect 31710 33690 31740 33810
rect 31860 33690 32700 33810
rect 32820 33690 32850 33810
rect 31710 33675 32850 33690
rect 31710 33660 31890 33675
rect 32670 33660 32850 33675
rect 33630 33825 33810 33840
rect 36510 33825 36690 33840
rect 33630 33810 36690 33825
rect 33630 33690 33660 33810
rect 33780 33690 36540 33810
rect 36660 33690 36690 33810
rect 33630 33675 36690 33690
rect 33630 33660 33810 33675
rect 36510 33660 36690 33675
rect 41790 33825 41970 33840
rect 43710 33825 43890 33840
rect 41790 33810 43890 33825
rect 41790 33690 41820 33810
rect 41940 33690 43740 33810
rect 43860 33690 43890 33810
rect 41790 33675 43890 33690
rect 41790 33660 41970 33675
rect 43710 33660 43890 33675
rect 47310 33825 47490 33840
rect 48030 33825 48210 33840
rect 47310 33810 48210 33825
rect 47310 33690 47340 33810
rect 47460 33690 48060 33810
rect 48180 33690 48210 33810
rect 47310 33675 48210 33690
rect 47310 33660 47490 33675
rect 48030 33660 48210 33675
rect 16830 33525 17010 33540
rect 17550 33525 17730 33540
rect 26670 33525 26850 33540
rect 16830 33510 26850 33525
rect 16830 33390 16860 33510
rect 16980 33390 17580 33510
rect 17700 33390 26700 33510
rect 26820 33390 26850 33510
rect 16830 33375 26850 33390
rect 16830 33360 17010 33375
rect 17550 33360 17730 33375
rect 26670 33360 26850 33375
rect 30990 33525 31170 33540
rect 31710 33525 31890 33540
rect 30990 33510 31890 33525
rect 30990 33390 31020 33510
rect 31140 33390 31740 33510
rect 31860 33390 31890 33510
rect 30990 33375 31890 33390
rect 30990 33360 31170 33375
rect 31710 33360 31890 33375
rect 37230 33525 37410 33540
rect 39390 33525 39570 33540
rect 37230 33510 39570 33525
rect 37230 33390 37260 33510
rect 37380 33390 39420 33510
rect 39540 33390 39570 33510
rect 37230 33375 39570 33390
rect 37230 33360 37410 33375
rect 39390 33360 39570 33375
rect 40110 33525 40290 33540
rect 40830 33525 41010 33540
rect 40110 33510 41010 33525
rect 40110 33390 40140 33510
rect 40260 33390 40860 33510
rect 40980 33390 41010 33510
rect 40110 33375 41010 33390
rect 40110 33360 40290 33375
rect 40830 33360 41010 33375
rect 41310 33525 41490 33540
rect 42270 33525 42450 33540
rect 41310 33510 42450 33525
rect 41310 33390 41340 33510
rect 41460 33390 42300 33510
rect 42420 33390 42450 33510
rect 41310 33375 42450 33390
rect 41310 33360 41490 33375
rect 42270 33360 42450 33375
rect 46110 33525 46290 33540
rect 46590 33525 46770 33540
rect 47550 33525 47730 33540
rect 46110 33510 47730 33525
rect 46110 33390 46140 33510
rect 46260 33390 46620 33510
rect 46740 33390 47580 33510
rect 47700 33390 47730 33510
rect 46110 33375 47730 33390
rect 46110 33360 46290 33375
rect 46590 33360 46770 33375
rect 47550 33360 47730 33375
rect 13470 33225 13650 33240
rect 13950 33225 14130 33240
rect 13470 33210 14130 33225
rect 13470 33090 13500 33210
rect 13620 33090 13980 33210
rect 14100 33090 14130 33210
rect 13470 33075 14130 33090
rect 13470 33060 13650 33075
rect 13950 33060 14130 33075
rect 15150 33225 15330 33240
rect 15870 33225 16050 33240
rect 16590 33225 16770 33240
rect 15150 33210 16770 33225
rect 15150 33090 15180 33210
rect 15300 33090 15900 33210
rect 16020 33090 16620 33210
rect 16740 33090 16770 33210
rect 15150 33075 16770 33090
rect 15150 33060 15330 33075
rect 15870 33060 16050 33075
rect 16590 33060 16770 33075
rect 18990 33225 19170 33240
rect 23790 33225 23970 33240
rect 18990 33210 23970 33225
rect 18990 33090 19020 33210
rect 19140 33090 23820 33210
rect 23940 33090 23970 33210
rect 18990 33075 23970 33090
rect 18990 33060 19170 33075
rect 23790 33060 23970 33075
rect 24750 33225 24930 33240
rect 25710 33225 25890 33240
rect 24750 33210 25890 33225
rect 24750 33090 24780 33210
rect 24900 33090 25740 33210
rect 25860 33090 25890 33210
rect 24750 33075 25890 33090
rect 24750 33060 24930 33075
rect 25710 33060 25890 33075
rect 33150 33225 33330 33240
rect 35070 33225 35250 33240
rect 33150 33210 35250 33225
rect 33150 33090 33180 33210
rect 33300 33090 35100 33210
rect 35220 33090 35250 33210
rect 33150 33075 35250 33090
rect 33150 33060 33330 33075
rect 35070 33060 35250 33075
rect 35790 33225 35970 33240
rect 39390 33225 39570 33240
rect 41070 33225 41250 33240
rect 42030 33225 42210 33240
rect 35790 33210 42210 33225
rect 35790 33090 35820 33210
rect 35940 33090 39420 33210
rect 39540 33090 41100 33210
rect 41220 33090 42060 33210
rect 42180 33090 42210 33210
rect 35790 33075 42210 33090
rect 35790 33060 35970 33075
rect 39390 33060 39570 33075
rect 41070 33060 41250 33075
rect 42030 33060 42210 33075
rect 43950 33225 44130 33240
rect 46590 33225 46770 33240
rect 43950 33210 46770 33225
rect 43950 33090 43980 33210
rect 44100 33090 46620 33210
rect 46740 33090 46770 33210
rect 43950 33075 46770 33090
rect 43950 33060 44130 33075
rect 46590 33060 46770 33075
rect 11550 32925 11730 32940
rect 15630 32925 15810 32940
rect 19470 32925 19650 32940
rect 11550 32910 19650 32925
rect 11550 32790 11580 32910
rect 11700 32790 15660 32910
rect 15780 32790 19500 32910
rect 19620 32790 19650 32910
rect 6510 32775 6690 32790
rect 0 32760 6690 32775
rect 11550 32775 19650 32790
rect 11550 32760 11730 32775
rect 15630 32760 15810 32775
rect 19470 32760 19650 32775
rect 21150 32925 21330 32940
rect 25230 32925 25410 32940
rect 21150 32910 25410 32925
rect 21150 32790 21180 32910
rect 21300 32790 25260 32910
rect 25380 32790 25410 32910
rect 21150 32775 25410 32790
rect 21150 32760 21330 32775
rect 25230 32760 25410 32775
rect 29070 32925 29250 32940
rect 34590 32925 34770 32940
rect 38190 32925 38370 32940
rect 29070 32910 38370 32925
rect 29070 32790 29100 32910
rect 29220 32790 34620 32910
rect 34740 32790 38220 32910
rect 38340 32790 38370 32910
rect 29070 32775 38370 32790
rect 29070 32760 29250 32775
rect 34590 32760 34770 32775
rect 38190 32760 38370 32775
rect 39870 32925 40050 32940
rect 45870 32925 46050 32940
rect 48030 32925 48210 32940
rect 39870 32910 48210 32925
rect 39870 32790 39900 32910
rect 40020 32790 45900 32910
rect 46020 32790 48060 32910
rect 48180 32790 48210 32910
rect 39870 32775 48210 32790
rect 39870 32760 40050 32775
rect 45870 32760 46050 32775
rect 48030 32760 48210 32775
rect 0 32640 6540 32760
rect 6660 32640 6690 32760
rect 0 32625 6690 32640
rect 6510 32610 6690 32625
rect 16350 32625 16530 32640
rect 17070 32625 17250 32640
rect 16350 32610 17250 32625
rect 16350 32490 16380 32610
rect 16500 32490 17100 32610
rect 17220 32490 17250 32610
rect 16350 32475 17250 32490
rect 16350 32460 16530 32475
rect 17070 32460 17250 32475
rect 36990 32625 37170 32640
rect 39630 32625 39810 32640
rect 36990 32610 39810 32625
rect 36990 32490 37020 32610
rect 37140 32490 39660 32610
rect 39780 32490 39810 32610
rect 36990 32475 39810 32490
rect 36990 32460 37170 32475
rect 39630 32460 39810 32475
rect 41310 32625 41490 32640
rect 50910 32625 51090 32640
rect 41310 32610 51090 32625
rect 41310 32490 41340 32610
rect 41460 32490 50940 32610
rect 51060 32490 51090 32610
rect 41310 32475 51090 32490
rect 41310 32460 41490 32475
rect 50910 32460 51090 32475
rect 10830 32325 11010 32340
rect 11790 32325 11970 32340
rect 10830 32310 11970 32325
rect 10830 32190 10860 32310
rect 10980 32190 11820 32310
rect 11940 32190 11970 32310
rect 10830 32175 11970 32190
rect 10830 32160 11010 32175
rect 11790 32160 11970 32175
rect 21630 32325 21810 32340
rect 26190 32325 26370 32340
rect 21630 32310 26370 32325
rect 21630 32190 21660 32310
rect 21780 32190 26220 32310
rect 26340 32190 26370 32310
rect 21630 32175 26370 32190
rect 21630 32160 21810 32175
rect 26190 32160 26370 32175
rect 41310 32025 41490 32040
rect 43950 32025 44130 32040
rect 44430 32025 44610 32040
rect 41310 32010 44610 32025
rect 41310 31890 41340 32010
rect 41460 31890 43980 32010
rect 44100 31890 44460 32010
rect 44580 31890 44610 32010
rect 41310 31875 44610 31890
rect 41310 31860 41490 31875
rect 43950 31860 44130 31875
rect 44430 31860 44610 31875
rect 6030 31725 6210 31740
rect 6990 31725 7170 31740
rect 6030 31710 7170 31725
rect 6030 31590 6060 31710
rect 6180 31590 7020 31710
rect 7140 31590 7170 31710
rect 6030 31575 7170 31590
rect 6030 31560 6210 31575
rect 6990 31560 7170 31575
rect 16830 31725 17010 31740
rect 17310 31725 17490 31740
rect 16830 31710 17490 31725
rect 16830 31590 16860 31710
rect 16980 31590 17340 31710
rect 17460 31590 17490 31710
rect 16830 31575 17490 31590
rect 16830 31560 17010 31575
rect 17310 31560 17490 31575
rect 35070 31725 35250 31740
rect 39390 31725 39570 31740
rect 35070 31710 39570 31725
rect 35070 31590 35100 31710
rect 35220 31590 39420 31710
rect 39540 31590 39570 31710
rect 35070 31575 39570 31590
rect 35070 31560 35250 31575
rect 39390 31560 39570 31575
rect 6270 31425 6450 31440
rect 8190 31425 8370 31440
rect 6270 31410 8370 31425
rect 6270 31290 6300 31410
rect 6420 31290 8220 31410
rect 8340 31290 8370 31410
rect 6270 31275 8370 31290
rect 6270 31260 6450 31275
rect 8190 31260 8370 31275
rect 19230 31425 19410 31440
rect 21150 31425 21330 31440
rect 22830 31425 23010 31440
rect 19230 31410 23010 31425
rect 19230 31290 19260 31410
rect 19380 31290 21180 31410
rect 21300 31290 22860 31410
rect 22980 31290 23010 31410
rect 19230 31275 23010 31290
rect 19230 31260 19410 31275
rect 21150 31260 21330 31275
rect 22830 31260 23010 31275
rect 25470 31425 25650 31440
rect 26910 31425 27090 31440
rect 25470 31410 27090 31425
rect 25470 31290 25500 31410
rect 25620 31290 26940 31410
rect 27060 31290 27090 31410
rect 25470 31275 27090 31290
rect 25470 31260 25650 31275
rect 26910 31260 27090 31275
rect 27390 31425 27570 31440
rect 29790 31425 29970 31440
rect 32190 31425 32370 31440
rect 35070 31425 35250 31440
rect 27390 31410 35250 31425
rect 27390 31290 27420 31410
rect 27540 31290 29820 31410
rect 29940 31290 32220 31410
rect 32340 31290 35100 31410
rect 35220 31290 35250 31410
rect 27390 31275 35250 31290
rect 27390 31260 27570 31275
rect 29790 31260 29970 31275
rect 32190 31260 32370 31275
rect 35070 31260 35250 31275
rect 43230 31425 43410 31440
rect 43950 31425 44130 31440
rect 45150 31425 45330 31440
rect 46590 31425 46770 31440
rect 43230 31410 46770 31425
rect 43230 31290 43260 31410
rect 43380 31290 43980 31410
rect 44100 31290 45180 31410
rect 45300 31290 46620 31410
rect 46740 31290 46770 31410
rect 43230 31275 46770 31290
rect 43230 31260 43410 31275
rect 43950 31260 44130 31275
rect 45150 31260 45330 31275
rect 46590 31260 46770 31275
rect 7950 31125 8130 31140
rect 9150 31125 9330 31140
rect 9630 31125 9810 31140
rect 7950 31110 9810 31125
rect 7950 30990 7980 31110
rect 8100 30990 9180 31110
rect 9300 30990 9660 31110
rect 9780 30990 9810 31110
rect 7950 30975 9810 30990
rect 7950 30960 8130 30975
rect 9150 30960 9330 30975
rect 9630 30960 9810 30975
rect 20910 31125 21090 31140
rect 21630 31125 21810 31140
rect 22590 31125 22770 31140
rect 24030 31125 24210 31140
rect 20910 31110 24210 31125
rect 20910 30990 20940 31110
rect 21060 30990 21660 31110
rect 21780 30990 22620 31110
rect 22740 30990 24060 31110
rect 24180 30990 24210 31110
rect 20910 30975 24210 30990
rect 20910 30960 21090 30975
rect 21630 30960 21810 30975
rect 22590 30960 22770 30975
rect 24030 30960 24210 30975
rect 25950 31125 26130 31140
rect 29070 31125 29250 31140
rect 25950 31110 29250 31125
rect 25950 30990 25980 31110
rect 26100 30990 29100 31110
rect 29220 30990 29250 31110
rect 25950 30975 29250 30990
rect 25950 30960 26130 30975
rect 29070 30960 29250 30975
rect 36750 31125 36930 31140
rect 38190 31125 38370 31140
rect 40830 31125 41010 31140
rect 36750 31110 41010 31125
rect 36750 30990 36780 31110
rect 36900 30990 38220 31110
rect 38340 30990 40860 31110
rect 40980 30990 41010 31110
rect 36750 30975 41010 30990
rect 36750 30960 36930 30975
rect 38190 30960 38370 30975
rect 40830 30960 41010 30975
rect 42750 31125 42930 31140
rect 43470 31125 43650 31140
rect 42750 31110 43650 31125
rect 42750 30990 42780 31110
rect 42900 30990 43500 31110
rect 43620 30990 43650 31110
rect 42750 30975 43650 30990
rect 42750 30960 42930 30975
rect 43470 30960 43650 30975
rect 8190 30825 8370 30840
rect 10110 30825 10290 30840
rect 13710 30825 13890 30840
rect 8190 30810 13890 30825
rect 8190 30690 8220 30810
rect 8340 30690 10140 30810
rect 10260 30690 13740 30810
rect 13860 30690 13890 30810
rect 8190 30675 13890 30690
rect 8190 30660 8370 30675
rect 10110 30660 10290 30675
rect 13710 30660 13890 30675
rect 18990 30825 19170 30840
rect 19950 30825 20130 30840
rect 18990 30810 20130 30825
rect 18990 30690 19020 30810
rect 19140 30690 19980 30810
rect 20100 30690 20130 30810
rect 18990 30675 20130 30690
rect 18990 30660 19170 30675
rect 19950 30660 20130 30675
rect 25710 30825 25890 30840
rect 27150 30825 27330 30840
rect 25710 30810 27330 30825
rect 25710 30690 25740 30810
rect 25860 30690 27180 30810
rect 27300 30690 27330 30810
rect 25710 30675 27330 30690
rect 25710 30660 25890 30675
rect 27150 30660 27330 30675
rect 29070 30825 29250 30840
rect 29550 30825 29730 30840
rect 29070 30810 29730 30825
rect 29070 30690 29100 30810
rect 29220 30690 29580 30810
rect 29700 30690 29730 30810
rect 29070 30675 29730 30690
rect 29070 30660 29250 30675
rect 29550 30660 29730 30675
rect 36270 30825 36450 30840
rect 36750 30825 36930 30840
rect 36270 30810 36930 30825
rect 36270 30690 36300 30810
rect 36420 30690 36780 30810
rect 36900 30690 36930 30810
rect 36270 30675 36930 30690
rect 36270 30660 36450 30675
rect 36750 30660 36930 30675
rect 39150 30825 39330 30840
rect 39630 30825 39810 30840
rect 39150 30810 39810 30825
rect 39150 30690 39180 30810
rect 39300 30690 39660 30810
rect 39780 30690 39810 30810
rect 39150 30675 39810 30690
rect 39150 30660 39330 30675
rect 39630 30660 39810 30675
rect 41550 30825 41730 30840
rect 43710 30825 43890 30840
rect 41550 30810 43890 30825
rect 41550 30690 41580 30810
rect 41700 30690 43740 30810
rect 43860 30690 43890 30810
rect 41550 30675 43890 30690
rect 41550 30660 41730 30675
rect 43710 30660 43890 30675
rect 44670 30825 44850 30840
rect 46110 30825 46290 30840
rect 44670 30810 46290 30825
rect 44670 30690 44700 30810
rect 44820 30690 46140 30810
rect 46260 30690 46290 30810
rect 44670 30675 46290 30690
rect 44670 30660 44850 30675
rect 46110 30660 46290 30675
rect 5310 30525 5490 30540
rect 8430 30525 8610 30540
rect 5310 30510 8610 30525
rect 5310 30390 5340 30510
rect 5460 30390 8460 30510
rect 8580 30390 8610 30510
rect 5310 30375 8610 30390
rect 5310 30360 5490 30375
rect 8430 30360 8610 30375
rect 11790 30525 11970 30540
rect 12990 30525 13170 30540
rect 11790 30510 13170 30525
rect 11790 30390 11820 30510
rect 11940 30390 13020 30510
rect 13140 30390 13170 30510
rect 11790 30375 13170 30390
rect 11790 30360 11970 30375
rect 12990 30360 13170 30375
rect 21150 30525 21330 30540
rect 21870 30525 22050 30540
rect 21150 30510 22050 30525
rect 21150 30390 21180 30510
rect 21300 30390 21900 30510
rect 22020 30390 22050 30510
rect 21150 30375 22050 30390
rect 21150 30360 21330 30375
rect 21870 30360 22050 30375
rect 26670 30525 26850 30540
rect 27390 30525 27570 30540
rect 28590 30525 28770 30540
rect 26670 30510 28770 30525
rect 26670 30390 26700 30510
rect 26820 30390 27420 30510
rect 27540 30390 28620 30510
rect 28740 30390 28770 30510
rect 26670 30375 28770 30390
rect 26670 30360 26850 30375
rect 27390 30360 27570 30375
rect 28590 30360 28770 30375
rect 33630 30525 33810 30540
rect 35070 30525 35250 30540
rect 33630 30510 35250 30525
rect 33630 30390 33660 30510
rect 33780 30390 35100 30510
rect 35220 30390 35250 30510
rect 33630 30375 35250 30390
rect 33630 30360 33810 30375
rect 35070 30360 35250 30375
rect 36030 30525 36210 30540
rect 37710 30525 37890 30540
rect 36030 30510 37890 30525
rect 36030 30390 36060 30510
rect 36180 30390 37740 30510
rect 37860 30390 37890 30510
rect 36030 30375 37890 30390
rect 36030 30360 36210 30375
rect 37710 30360 37890 30375
rect 40350 30525 40530 30540
rect 44910 30525 45090 30540
rect 40350 30510 45090 30525
rect 40350 30390 40380 30510
rect 40500 30390 44940 30510
rect 45060 30390 45090 30510
rect 40350 30375 45090 30390
rect 40350 30360 40530 30375
rect 44910 30360 45090 30375
rect 9390 30225 9570 30240
rect 12030 30225 12210 30240
rect 9390 30210 12210 30225
rect 9390 30090 9420 30210
rect 9540 30090 12060 30210
rect 12180 30090 12210 30210
rect 9390 30075 12210 30090
rect 9390 30060 9570 30075
rect 12030 30060 12210 30075
rect 17070 30225 17250 30240
rect 17550 30225 17730 30240
rect 20910 30225 21090 30240
rect 17070 30210 21090 30225
rect 17070 30090 17100 30210
rect 17220 30090 17580 30210
rect 17700 30090 20940 30210
rect 21060 30090 21090 30210
rect 17070 30075 21090 30090
rect 17070 30060 17250 30075
rect 17550 30060 17730 30075
rect 20910 30060 21090 30075
rect 28590 30225 28770 30240
rect 30030 30225 30210 30240
rect 28590 30210 30210 30225
rect 28590 30090 28620 30210
rect 28740 30090 30060 30210
rect 30180 30090 30210 30210
rect 28590 30075 30210 30090
rect 28590 30060 28770 30075
rect 30030 30060 30210 30075
rect 35070 30225 35250 30240
rect 35550 30225 35730 30240
rect 35070 30210 35730 30225
rect 35070 30090 35100 30210
rect 35220 30090 35580 30210
rect 35700 30090 35730 30210
rect 35070 30075 35730 30090
rect 35070 30060 35250 30075
rect 35550 30060 35730 30075
rect 43710 30225 43890 30240
rect 47550 30225 47730 30240
rect 43710 30210 47730 30225
rect 43710 30090 43740 30210
rect 43860 30090 47580 30210
rect 47700 30090 47730 30210
rect 43710 30075 47730 30090
rect 43710 30060 43890 30075
rect 47550 30060 47730 30075
rect 12030 29925 12210 29940
rect 22110 29925 22290 29940
rect 12030 29910 22290 29925
rect 12030 29790 12060 29910
rect 12180 29790 22140 29910
rect 22260 29790 22290 29910
rect 12030 29775 22290 29790
rect 12030 29760 12210 29775
rect 22110 29760 22290 29775
rect 28350 29925 28530 29940
rect 29070 29925 29250 29940
rect 28350 29910 29250 29925
rect 28350 29790 28380 29910
rect 28500 29790 29100 29910
rect 29220 29790 29250 29910
rect 28350 29775 29250 29790
rect 28350 29760 28530 29775
rect 29070 29760 29250 29775
rect 34830 29925 35010 29940
rect 35550 29925 35730 29940
rect 34830 29910 35730 29925
rect 34830 29790 34860 29910
rect 34980 29790 35580 29910
rect 35700 29790 35730 29910
rect 34830 29775 35730 29790
rect 34830 29760 35010 29775
rect 35550 29760 35730 29775
rect 38430 29925 38610 29940
rect 43950 29925 44130 29940
rect 38430 29910 44130 29925
rect 38430 29790 38460 29910
rect 38580 29790 43980 29910
rect 44100 29790 44130 29910
rect 38430 29775 44130 29790
rect 38430 29760 38610 29775
rect 43950 29760 44130 29775
rect 9150 29625 9330 29640
rect 9870 29625 10050 29640
rect 9150 29610 10050 29625
rect 9150 29490 9180 29610
rect 9300 29490 9900 29610
rect 10020 29490 10050 29610
rect 9150 29475 10050 29490
rect 9150 29460 9330 29475
rect 9870 29460 10050 29475
rect 17790 29625 17970 29640
rect 19710 29625 19890 29640
rect 17790 29610 19890 29625
rect 17790 29490 17820 29610
rect 17940 29490 19740 29610
rect 19860 29490 19890 29610
rect 17790 29475 19890 29490
rect 17790 29460 17970 29475
rect 19710 29460 19890 29475
rect 25470 29625 25650 29640
rect 27630 29625 27810 29640
rect 33870 29625 34050 29640
rect 25470 29610 34050 29625
rect 25470 29490 25500 29610
rect 25620 29490 27660 29610
rect 27780 29490 33900 29610
rect 34020 29490 34050 29610
rect 25470 29475 34050 29490
rect 25470 29460 25650 29475
rect 27630 29460 27810 29475
rect 33870 29460 34050 29475
rect 26910 29325 27090 29340
rect 33630 29325 33810 29340
rect 26910 29310 33810 29325
rect 26910 29190 26940 29310
rect 27060 29190 33660 29310
rect 33780 29190 33810 29310
rect 26910 29175 33810 29190
rect 26910 29160 27090 29175
rect 33630 29160 33810 29175
rect 35070 28425 35250 28440
rect 37950 28425 38130 28440
rect 35070 28410 38130 28425
rect 35070 28290 35100 28410
rect 35220 28290 37980 28410
rect 38100 28290 38130 28410
rect 35070 28275 38130 28290
rect 35070 28260 35250 28275
rect 37950 28260 38130 28275
rect 12510 28125 12690 28140
rect 21630 28125 21810 28140
rect 12510 28110 21810 28125
rect 12510 27990 12540 28110
rect 12660 27990 21660 28110
rect 21780 27990 21810 28110
rect 12510 27975 21810 27990
rect 12510 27960 12690 27975
rect 21630 27960 21810 27975
rect 23070 28125 23250 28140
rect 23550 28125 23730 28140
rect 25470 28125 25650 28140
rect 23070 28110 25650 28125
rect 23070 27990 23100 28110
rect 23220 27990 23580 28110
rect 23700 27990 25500 28110
rect 25620 27990 25650 28110
rect 23070 27975 25650 27990
rect 23070 27960 23250 27975
rect 23550 27960 23730 27975
rect 25470 27960 25650 27975
rect 33150 28125 33330 28140
rect 35310 28125 35490 28140
rect 33150 28110 35490 28125
rect 33150 27990 33180 28110
rect 33300 27990 35340 28110
rect 35460 27990 35490 28110
rect 33150 27975 35490 27990
rect 33150 27960 33330 27975
rect 35310 27960 35490 27975
rect 36510 28125 36690 28140
rect 42030 28125 42210 28140
rect 43710 28125 43890 28140
rect 36510 28110 43890 28125
rect 36510 27990 36540 28110
rect 36660 27990 42060 28110
rect 42180 27990 43740 28110
rect 43860 27990 43890 28110
rect 36510 27975 43890 27990
rect 36510 27960 36690 27975
rect 42030 27960 42210 27975
rect 43710 27960 43890 27975
rect 11310 27825 11490 27840
rect 12750 27825 12930 27840
rect 13230 27825 13410 27840
rect 11310 27810 13410 27825
rect 11310 27690 11340 27810
rect 11460 27690 12780 27810
rect 12900 27690 13260 27810
rect 13380 27690 13410 27810
rect 11310 27675 13410 27690
rect 11310 27660 11490 27675
rect 12750 27660 12930 27675
rect 13230 27660 13410 27675
rect 15150 27825 15330 27840
rect 15870 27825 16050 27840
rect 15150 27810 16050 27825
rect 15150 27690 15180 27810
rect 15300 27690 15900 27810
rect 16020 27690 16050 27810
rect 15150 27675 16050 27690
rect 15150 27660 15330 27675
rect 15870 27660 16050 27675
rect 17790 27825 17970 27840
rect 21630 27825 21810 27840
rect 24030 27825 24210 27840
rect 32910 27825 33090 27840
rect 17790 27810 33090 27825
rect 17790 27690 17820 27810
rect 17940 27690 21660 27810
rect 21780 27690 24060 27810
rect 24180 27690 32940 27810
rect 33060 27690 33090 27810
rect 17790 27675 33090 27690
rect 17790 27660 17970 27675
rect 21630 27660 21810 27675
rect 24030 27660 24210 27675
rect 32910 27660 33090 27675
rect 38910 27825 39090 27840
rect 46590 27825 46770 27840
rect 38910 27810 46770 27825
rect 38910 27690 38940 27810
rect 39060 27690 46620 27810
rect 46740 27690 46770 27810
rect 38910 27675 46770 27690
rect 38910 27660 39090 27675
rect 46590 27660 46770 27675
rect 48750 27825 48930 27840
rect 49950 27825 50130 27840
rect 48750 27810 50130 27825
rect 48750 27690 48780 27810
rect 48900 27690 49980 27810
rect 50100 27690 50130 27810
rect 48750 27675 50130 27690
rect 48750 27660 48930 27675
rect 49950 27660 50130 27675
rect 7710 27510 7890 27540
rect 7710 27390 7740 27510
rect 7860 27390 7890 27510
rect 6030 27375 6210 27390
rect 0 27360 6210 27375
rect 7710 27360 7890 27390
rect 8670 27525 8850 27540
rect 9150 27525 9330 27540
rect 8670 27510 9330 27525
rect 8670 27390 8700 27510
rect 8820 27390 9180 27510
rect 9300 27390 9330 27510
rect 8670 27375 9330 27390
rect 8670 27360 8850 27375
rect 9150 27360 9330 27375
rect 13230 27525 13410 27540
rect 15390 27525 15570 27540
rect 13230 27510 15570 27525
rect 13230 27390 13260 27510
rect 13380 27390 15420 27510
rect 15540 27390 15570 27510
rect 13230 27375 15570 27390
rect 13230 27360 13410 27375
rect 15390 27360 15570 27375
rect 19230 27525 19410 27540
rect 23310 27525 23490 27540
rect 19230 27510 23490 27525
rect 19230 27390 19260 27510
rect 19380 27390 23340 27510
rect 23460 27390 23490 27510
rect 19230 27375 23490 27390
rect 19230 27360 19410 27375
rect 23310 27360 23490 27375
rect 24510 27525 24690 27540
rect 25470 27525 25650 27540
rect 24510 27510 25650 27525
rect 24510 27390 24540 27510
rect 24660 27390 25500 27510
rect 25620 27390 25650 27510
rect 24510 27375 25650 27390
rect 24510 27360 24690 27375
rect 25470 27360 25650 27375
rect 28350 27525 28530 27540
rect 28830 27525 29010 27540
rect 28350 27510 29010 27525
rect 28350 27390 28380 27510
rect 28500 27390 28860 27510
rect 28980 27390 29010 27510
rect 28350 27375 29010 27390
rect 28350 27360 28530 27375
rect 28830 27360 29010 27375
rect 30270 27525 30450 27540
rect 32190 27525 32370 27540
rect 30270 27510 32370 27525
rect 30270 27390 30300 27510
rect 30420 27390 32220 27510
rect 32340 27390 32370 27510
rect 30270 27375 32370 27390
rect 30270 27360 30450 27375
rect 32190 27360 32370 27375
rect 35790 27525 35970 27540
rect 38430 27525 38610 27540
rect 35790 27510 38610 27525
rect 35790 27390 35820 27510
rect 35940 27390 38460 27510
rect 38580 27390 38610 27510
rect 35790 27375 38610 27390
rect 35790 27360 35970 27375
rect 38430 27360 38610 27375
rect 48510 27525 48690 27540
rect 48990 27525 49170 27540
rect 48510 27510 49170 27525
rect 48510 27390 48540 27510
rect 48660 27390 49020 27510
rect 49140 27390 49170 27510
rect 48510 27375 49170 27390
rect 48510 27360 48690 27375
rect 48990 27360 49170 27375
rect 0 27240 6060 27360
rect 6180 27240 6210 27360
rect 0 27225 6210 27240
rect 6030 27210 6210 27225
rect 7725 26640 7875 27360
rect 11070 27225 11250 27240
rect 12510 27225 12690 27240
rect 11070 27210 12690 27225
rect 11070 27090 11100 27210
rect 11220 27090 12540 27210
rect 12660 27090 12690 27210
rect 11070 27075 12690 27090
rect 11070 27060 11250 27075
rect 12510 27060 12690 27075
rect 16590 27225 16770 27240
rect 18030 27225 18210 27240
rect 16590 27210 18210 27225
rect 16590 27090 16620 27210
rect 16740 27090 18060 27210
rect 18180 27090 18210 27210
rect 16590 27075 18210 27090
rect 16590 27060 16770 27075
rect 18030 27060 18210 27075
rect 20670 27225 20850 27240
rect 21150 27225 21330 27240
rect 25230 27225 25410 27240
rect 20670 27210 25410 27225
rect 20670 27090 20700 27210
rect 20820 27090 21180 27210
rect 21300 27090 25260 27210
rect 25380 27090 25410 27210
rect 20670 27075 25410 27090
rect 20670 27060 20850 27075
rect 21150 27060 21330 27075
rect 25230 27060 25410 27075
rect 31950 27225 32130 27240
rect 34350 27225 34530 27240
rect 31950 27210 34530 27225
rect 31950 27090 31980 27210
rect 32100 27090 34380 27210
rect 34500 27090 34530 27210
rect 31950 27075 34530 27090
rect 31950 27060 32130 27075
rect 34350 27060 34530 27075
rect 36030 27225 36210 27240
rect 36510 27225 36690 27240
rect 36030 27210 36690 27225
rect 36030 27090 36060 27210
rect 36180 27090 36540 27210
rect 36660 27090 36690 27210
rect 36030 27075 36690 27090
rect 36030 27060 36210 27075
rect 36510 27060 36690 27075
rect 38430 27225 38610 27240
rect 41310 27225 41490 27240
rect 43470 27225 43650 27240
rect 38430 27210 43650 27225
rect 38430 27090 38460 27210
rect 38580 27090 41340 27210
rect 41460 27090 43500 27210
rect 43620 27090 43650 27210
rect 38430 27075 43650 27090
rect 38430 27060 38610 27075
rect 41310 27060 41490 27075
rect 43470 27060 43650 27075
rect 46830 27225 47010 27240
rect 48030 27225 48210 27240
rect 46830 27210 48210 27225
rect 46830 27090 46860 27210
rect 46980 27090 48060 27210
rect 48180 27090 48210 27210
rect 46830 27075 48210 27090
rect 46830 27060 47010 27075
rect 48030 27060 48210 27075
rect 8670 26925 8850 26940
rect 10350 26925 10530 26940
rect 18750 26925 18930 26940
rect 8670 26910 18930 26925
rect 8670 26790 8700 26910
rect 8820 26790 10380 26910
rect 10500 26790 18780 26910
rect 18900 26790 18930 26910
rect 8670 26775 18930 26790
rect 8670 26760 8850 26775
rect 10350 26760 10530 26775
rect 18750 26760 18930 26775
rect 30750 26925 30930 26940
rect 32430 26925 32610 26940
rect 30750 26910 32610 26925
rect 30750 26790 30780 26910
rect 30900 26790 32460 26910
rect 32580 26790 32610 26910
rect 30750 26775 32610 26790
rect 30750 26760 30930 26775
rect 32430 26760 32610 26775
rect 36510 26925 36690 26940
rect 38670 26925 38850 26940
rect 36510 26910 38850 26925
rect 36510 26790 36540 26910
rect 36660 26790 38700 26910
rect 38820 26790 38850 26910
rect 36510 26775 38850 26790
rect 36510 26760 36690 26775
rect 38670 26760 38850 26775
rect 46830 26925 47010 26940
rect 48990 26925 49170 26940
rect 46830 26910 49170 26925
rect 46830 26790 46860 26910
rect 46980 26790 49020 26910
rect 49140 26790 49170 26910
rect 46830 26775 49170 26790
rect 46830 26760 47010 26775
rect 48990 26760 49170 26775
rect 7710 26610 7890 26640
rect 7710 26490 7740 26610
rect 7860 26490 7890 26610
rect 7710 26460 7890 26490
rect 15150 26625 15330 26640
rect 24030 26625 24210 26640
rect 15150 26610 24210 26625
rect 15150 26490 15180 26610
rect 15300 26490 24060 26610
rect 24180 26490 24210 26610
rect 15150 26475 24210 26490
rect 15150 26460 15330 26475
rect 24030 26460 24210 26475
rect 25710 26625 25890 26640
rect 36030 26625 36210 26640
rect 25710 26610 36210 26625
rect 25710 26490 25740 26610
rect 25860 26490 36060 26610
rect 36180 26490 36210 26610
rect 25710 26475 36210 26490
rect 25710 26460 25890 26475
rect 36030 26460 36210 26475
rect 43470 26625 43650 26640
rect 46590 26625 46770 26640
rect 43470 26610 46770 26625
rect 43470 26490 43500 26610
rect 43620 26490 46620 26610
rect 46740 26490 46770 26610
rect 43470 26475 46770 26490
rect 43470 26460 43650 26475
rect 46590 26460 46770 26475
rect 750 26325 930 26340
rect 15390 26325 15570 26340
rect 34590 26325 34770 26340
rect 750 26310 34770 26325
rect 750 26190 780 26310
rect 900 26190 15420 26310
rect 15540 26190 34620 26310
rect 34740 26190 34770 26310
rect 750 26175 34770 26190
rect 750 26160 930 26175
rect 15390 26160 15570 26175
rect 34590 26160 34770 26175
rect 9390 26025 9570 26040
rect 10110 26025 10290 26040
rect 9390 26010 10290 26025
rect 9390 25890 9420 26010
rect 9540 25890 10140 26010
rect 10260 25890 10290 26010
rect 9390 25875 10290 25890
rect 9390 25860 9570 25875
rect 10110 25860 10290 25875
rect 17070 26025 17250 26040
rect 17550 26025 17730 26040
rect 17070 26010 17730 26025
rect 17070 25890 17100 26010
rect 17220 25890 17580 26010
rect 17700 25890 17730 26010
rect 17070 25875 17730 25890
rect 17070 25860 17250 25875
rect 17550 25860 17730 25875
rect 25470 26025 25650 26040
rect 35550 26025 35730 26040
rect 25470 26010 35730 26025
rect 25470 25890 25500 26010
rect 25620 25890 35580 26010
rect 35700 25890 35730 26010
rect 25470 25875 35730 25890
rect 25470 25860 25650 25875
rect 35550 25860 35730 25875
rect 39150 25725 39330 25740
rect 42510 25725 42690 25740
rect 45870 25725 46050 25740
rect 39150 25710 46050 25725
rect 39150 25590 39180 25710
rect 39300 25590 42540 25710
rect 42660 25590 45900 25710
rect 46020 25590 46050 25710
rect 39150 25575 46050 25590
rect 39150 25560 39330 25575
rect 42510 25560 42690 25575
rect 45870 25560 46050 25575
rect 8430 25425 8610 25440
rect 9390 25425 9570 25440
rect 8430 25410 9570 25425
rect 8430 25290 8460 25410
rect 8580 25290 9420 25410
rect 9540 25290 9570 25410
rect 8430 25275 9570 25290
rect 8430 25260 8610 25275
rect 9390 25260 9570 25275
rect 12030 25425 12210 25440
rect 12990 25425 13170 25440
rect 12030 25410 13170 25425
rect 12030 25290 12060 25410
rect 12180 25290 13020 25410
rect 13140 25290 13170 25410
rect 12030 25275 13170 25290
rect 12030 25260 12210 25275
rect 12990 25260 13170 25275
rect 30510 25425 30690 25440
rect 31710 25425 31890 25440
rect 32670 25425 32850 25440
rect 30510 25410 32850 25425
rect 30510 25290 30540 25410
rect 30660 25290 31740 25410
rect 31860 25290 32700 25410
rect 32820 25290 32850 25410
rect 30510 25275 32850 25290
rect 30510 25260 30690 25275
rect 31710 25260 31890 25275
rect 32670 25260 32850 25275
rect 38670 25425 38850 25440
rect 39150 25425 39330 25440
rect 38670 25410 39330 25425
rect 38670 25290 38700 25410
rect 38820 25290 39180 25410
rect 39300 25290 39330 25410
rect 38670 25275 39330 25290
rect 38670 25260 38850 25275
rect 39150 25260 39330 25275
rect 40110 25425 40290 25440
rect 41070 25425 41250 25440
rect 43710 25425 43890 25440
rect 46110 25425 46290 25440
rect 40110 25410 46290 25425
rect 40110 25290 40140 25410
rect 40260 25290 41100 25410
rect 41220 25290 43740 25410
rect 43860 25290 46140 25410
rect 46260 25290 46290 25410
rect 40110 25275 46290 25290
rect 40110 25260 40290 25275
rect 41070 25260 41250 25275
rect 43710 25260 43890 25275
rect 46110 25260 46290 25275
rect 5310 25125 5490 25140
rect 6990 25125 7170 25140
rect 5310 25110 7170 25125
rect 5310 24990 5340 25110
rect 5460 24990 7020 25110
rect 7140 24990 7170 25110
rect 5310 24975 7170 24990
rect 5310 24960 5490 24975
rect 6990 24960 7170 24975
rect 8670 25125 8850 25140
rect 10830 25125 11010 25140
rect 8670 25110 11010 25125
rect 8670 24990 8700 25110
rect 8820 24990 10860 25110
rect 10980 24990 11010 25110
rect 8670 24975 11010 24990
rect 8670 24960 8850 24975
rect 10830 24960 11010 24975
rect 13470 25125 13650 25140
rect 14190 25125 14370 25140
rect 15390 25125 15570 25140
rect 13470 25110 15570 25125
rect 13470 24990 13500 25110
rect 13620 24990 14220 25110
rect 14340 24990 15420 25110
rect 15540 24990 15570 25110
rect 13470 24975 15570 24990
rect 13470 24960 13650 24975
rect 14190 24960 14370 24975
rect 15390 24960 15570 24975
rect 22350 25125 22530 25140
rect 24270 25125 24450 25140
rect 22350 25110 24450 25125
rect 22350 24990 22380 25110
rect 22500 24990 24300 25110
rect 24420 24990 24450 25110
rect 22350 24975 24450 24990
rect 22350 24960 22530 24975
rect 24270 24960 24450 24975
rect 27870 25125 28050 25140
rect 30510 25125 30690 25140
rect 27870 25110 30690 25125
rect 27870 24990 27900 25110
rect 28020 24990 30540 25110
rect 30660 24990 30690 25110
rect 27870 24975 30690 24990
rect 27870 24960 28050 24975
rect 30510 24960 30690 24975
rect 33150 25125 33330 25140
rect 35550 25125 35730 25140
rect 38910 25125 39090 25140
rect 39390 25125 39570 25140
rect 33150 25110 39570 25125
rect 33150 24990 33180 25110
rect 33300 24990 35580 25110
rect 35700 24990 38940 25110
rect 39060 24990 39420 25110
rect 39540 24990 39570 25110
rect 33150 24975 39570 24990
rect 33150 24960 33330 24975
rect 35550 24960 35730 24975
rect 38910 24960 39090 24975
rect 39390 24960 39570 24975
rect 40350 25125 40530 25140
rect 40830 25125 41010 25140
rect 40350 25110 41010 25125
rect 40350 24990 40380 25110
rect 40500 24990 40860 25110
rect 40980 24990 41010 25110
rect 40350 24975 41010 24990
rect 40350 24960 40530 24975
rect 40830 24960 41010 24975
rect 44430 25125 44610 25140
rect 47310 25125 47490 25140
rect 44430 25110 47490 25125
rect 44430 24990 44460 25110
rect 44580 24990 47340 25110
rect 47460 24990 47490 25110
rect 44430 24975 47490 24990
rect 44430 24960 44610 24975
rect 47310 24960 47490 24975
rect 6750 24825 6930 24840
rect 10110 24825 10290 24840
rect 6750 24810 10290 24825
rect 6750 24690 6780 24810
rect 6900 24690 10140 24810
rect 10260 24690 10290 24810
rect 6750 24675 10290 24690
rect 6750 24660 6930 24675
rect 10110 24660 10290 24675
rect 13470 24825 13650 24840
rect 15630 24825 15810 24840
rect 13470 24810 15810 24825
rect 13470 24690 13500 24810
rect 13620 24690 15660 24810
rect 15780 24690 15810 24810
rect 13470 24675 15810 24690
rect 13470 24660 13650 24675
rect 15630 24660 15810 24675
rect 27150 24825 27330 24840
rect 29310 24825 29490 24840
rect 27150 24810 29490 24825
rect 27150 24690 27180 24810
rect 27300 24690 29340 24810
rect 29460 24690 29490 24810
rect 27150 24675 29490 24690
rect 27150 24660 27330 24675
rect 29310 24660 29490 24675
rect 35790 24825 35970 24840
rect 35790 24810 41475 24825
rect 35790 24690 35820 24810
rect 35940 24690 41475 24810
rect 35790 24675 41475 24690
rect 55200 24675 55350 24690
rect 35790 24660 35970 24675
rect 7470 24525 7650 24540
rect 8670 24525 8850 24540
rect 7470 24510 8850 24525
rect 7470 24390 7500 24510
rect 7620 24390 8700 24510
rect 8820 24390 8850 24510
rect 7470 24375 8850 24390
rect 7470 24360 7650 24375
rect 8670 24360 8850 24375
rect 23070 24525 23250 24540
rect 23550 24525 23730 24540
rect 23070 24510 23730 24525
rect 23070 24390 23100 24510
rect 23220 24390 23580 24510
rect 23700 24390 23730 24510
rect 23070 24375 23730 24390
rect 23070 24360 23250 24375
rect 23550 24360 23730 24375
rect 29310 24525 29490 24540
rect 33630 24525 33810 24540
rect 29310 24510 33810 24525
rect 29310 24390 29340 24510
rect 29460 24390 33660 24510
rect 33780 24390 33810 24510
rect 29310 24375 33810 24390
rect 29310 24360 29490 24375
rect 33630 24360 33810 24375
rect 35310 24525 35490 24540
rect 37950 24525 38130 24540
rect 40830 24525 41010 24540
rect 41325 24525 55350 24675
rect 35310 24510 41010 24525
rect 55200 24510 55350 24525
rect 35310 24390 35340 24510
rect 35460 24390 37980 24510
rect 38100 24390 40860 24510
rect 40980 24390 41010 24510
rect 35310 24375 41010 24390
rect 35310 24360 35490 24375
rect 37950 24360 38130 24375
rect 40830 24360 41010 24375
rect 30750 24225 30930 24240
rect 31710 24225 31890 24240
rect 30750 24210 31890 24225
rect 30750 24090 30780 24210
rect 30900 24090 31740 24210
rect 31860 24090 31890 24210
rect 30750 24075 31890 24090
rect 30750 24060 30930 24075
rect 31710 24060 31890 24075
rect 32910 24225 33090 24240
rect 33630 24225 33810 24240
rect 32910 24210 33810 24225
rect 32910 24090 32940 24210
rect 33060 24090 33660 24210
rect 33780 24090 33810 24210
rect 32910 24075 33810 24090
rect 32910 24060 33090 24075
rect 33630 24060 33810 24075
rect 39630 24225 39810 24240
rect 42270 24225 42450 24240
rect 39630 24210 42450 24225
rect 39630 24090 39660 24210
rect 39780 24090 42300 24210
rect 42420 24090 42450 24210
rect 39630 24075 42450 24090
rect 39630 24060 39810 24075
rect 42270 24060 42450 24075
rect 24510 23925 24690 23940
rect 35790 23925 35970 23940
rect 24510 23910 35970 23925
rect 24510 23790 24540 23910
rect 24660 23790 35820 23910
rect 35940 23790 35970 23910
rect 24510 23775 35970 23790
rect 24510 23760 24690 23775
rect 35790 23760 35970 23775
rect 36510 23925 36690 23940
rect 39390 23925 39570 23940
rect 36510 23910 39570 23925
rect 36510 23790 36540 23910
rect 36660 23790 39420 23910
rect 39540 23790 39570 23910
rect 36510 23775 39570 23790
rect 36510 23760 36690 23775
rect 39390 23760 39570 23775
rect 12030 23625 12210 23640
rect 13950 23625 14130 23640
rect 12030 23610 14130 23625
rect 12030 23490 12060 23610
rect 12180 23490 13980 23610
rect 14100 23490 14130 23610
rect 12030 23475 14130 23490
rect 12030 23460 12210 23475
rect 13950 23460 14130 23475
rect 19710 23625 19890 23640
rect 25470 23625 25650 23640
rect 19710 23610 25650 23625
rect 19710 23490 19740 23610
rect 19860 23490 25500 23610
rect 25620 23490 25650 23610
rect 19710 23475 25650 23490
rect 19710 23460 19890 23475
rect 25470 23460 25650 23475
rect 28110 23625 28290 23640
rect 29070 23625 29250 23640
rect 28110 23610 29250 23625
rect 28110 23490 28140 23610
rect 28260 23490 29100 23610
rect 29220 23490 29250 23610
rect 28110 23475 29250 23490
rect 28110 23460 28290 23475
rect 29070 23460 29250 23475
rect 35070 23625 35250 23640
rect 36270 23625 36450 23640
rect 35070 23610 36450 23625
rect 35070 23490 35100 23610
rect 35220 23490 36300 23610
rect 36420 23490 36450 23610
rect 35070 23475 36450 23490
rect 35070 23460 35250 23475
rect 36270 23460 36450 23475
rect 40590 23625 40770 23640
rect 47790 23625 47970 23640
rect 40590 23610 47970 23625
rect 40590 23490 40620 23610
rect 40740 23490 47820 23610
rect 47940 23490 47970 23610
rect 40590 23475 47970 23490
rect 40590 23460 40770 23475
rect 47790 23460 47970 23475
rect 18030 23025 18210 23040
rect 18510 23025 18690 23040
rect 18030 23010 18690 23025
rect 18030 22890 18060 23010
rect 18180 22890 18540 23010
rect 18660 22890 18690 23010
rect 18030 22875 18690 22890
rect 18030 22860 18210 22875
rect 18510 22860 18690 22875
rect 20190 23025 20370 23040
rect 21150 23025 21330 23040
rect 20190 23010 21330 23025
rect 20190 22890 20220 23010
rect 20340 22890 21180 23010
rect 21300 22890 21330 23010
rect 20190 22875 21330 22890
rect 20190 22860 20370 22875
rect 21150 22860 21330 22875
rect 14190 22725 14370 22740
rect 21150 22725 21330 22740
rect 14190 22710 21330 22725
rect 14190 22590 14220 22710
rect 14340 22590 21180 22710
rect 21300 22590 21330 22710
rect 14190 22575 21330 22590
rect 14190 22560 14370 22575
rect 21150 22560 21330 22575
rect 18030 22425 18210 22440
rect 19710 22425 19890 22440
rect 18030 22410 19890 22425
rect 18030 22290 18060 22410
rect 18180 22290 19740 22410
rect 19860 22290 19890 22410
rect 18030 22275 19890 22290
rect 18030 22260 18210 22275
rect 19710 22260 19890 22275
rect 36270 22425 36450 22440
rect 36990 22425 37170 22440
rect 36270 22410 37170 22425
rect 36270 22290 36300 22410
rect 36420 22290 37020 22410
rect 37140 22290 37170 22410
rect 36270 22275 37170 22290
rect 36270 22260 36450 22275
rect 36990 22260 37170 22275
rect 6030 22125 6210 22140
rect 5325 22110 6210 22125
rect 5325 21990 6060 22110
rect 6180 21990 6210 22110
rect 5325 21975 6210 21990
rect 0 21825 5475 21975
rect 6030 21960 6210 21975
rect 32670 22125 32850 22140
rect 48990 22125 49170 22140
rect 32670 22110 49170 22125
rect 32670 21990 32700 22110
rect 32820 21990 49020 22110
rect 49140 21990 49170 22110
rect 32670 21975 49170 21990
rect 32670 21960 32850 21975
rect 48990 21960 49170 21975
rect 9630 21825 9810 21840
rect 10350 21825 10530 21840
rect 9630 21810 10530 21825
rect 9630 21690 9660 21810
rect 9780 21690 10380 21810
rect 10500 21690 10530 21810
rect 9630 21675 10530 21690
rect 9630 21660 9810 21675
rect 10350 21660 10530 21675
rect 22590 21825 22770 21840
rect 25470 21825 25650 21840
rect 22590 21810 25650 21825
rect 22590 21690 22620 21810
rect 22740 21690 25500 21810
rect 25620 21690 25650 21810
rect 22590 21675 25650 21690
rect 22590 21660 22770 21675
rect 25470 21660 25650 21675
rect 27870 21825 28050 21840
rect 28830 21825 29010 21840
rect 27870 21810 29010 21825
rect 27870 21690 27900 21810
rect 28020 21690 28860 21810
rect 28980 21690 29010 21810
rect 27870 21675 29010 21690
rect 27870 21660 28050 21675
rect 28830 21660 29010 21675
rect 38910 21825 39090 21840
rect 39870 21825 40050 21840
rect 38910 21810 40050 21825
rect 38910 21690 38940 21810
rect 39060 21690 39900 21810
rect 40020 21690 40050 21810
rect 38910 21675 40050 21690
rect 38910 21660 39090 21675
rect 39870 21660 40050 21675
rect 42030 21825 42210 21840
rect 43950 21825 44130 21840
rect 42030 21810 44130 21825
rect 42030 21690 42060 21810
rect 42180 21690 43980 21810
rect 44100 21690 44130 21810
rect 42030 21675 44130 21690
rect 42030 21660 42210 21675
rect 43950 21660 44130 21675
rect 6990 21525 7170 21540
rect 10350 21525 10530 21540
rect 6990 21510 10530 21525
rect 6990 21390 7020 21510
rect 7140 21390 10380 21510
rect 10500 21390 10530 21510
rect 6990 21375 10530 21390
rect 6990 21360 7170 21375
rect 10350 21360 10530 21375
rect 22110 21525 22290 21540
rect 23070 21525 23250 21540
rect 22110 21510 23250 21525
rect 22110 21390 22140 21510
rect 22260 21390 23100 21510
rect 23220 21390 23250 21510
rect 22110 21375 23250 21390
rect 22110 21360 22290 21375
rect 23070 21360 23250 21375
rect 26190 21525 26370 21540
rect 26670 21525 26850 21540
rect 26190 21510 26850 21525
rect 26190 21390 26220 21510
rect 26340 21390 26700 21510
rect 26820 21390 26850 21510
rect 26190 21375 26850 21390
rect 26190 21360 26370 21375
rect 26670 21360 26850 21375
rect 36750 21525 36930 21540
rect 42030 21525 42210 21540
rect 43710 21525 43890 21540
rect 47310 21525 47490 21540
rect 48030 21525 48210 21540
rect 36750 21510 44835 21525
rect 36750 21390 36780 21510
rect 36900 21390 42060 21510
rect 42180 21390 43740 21510
rect 43860 21390 44835 21510
rect 36750 21375 44835 21390
rect 36750 21360 36930 21375
rect 42030 21360 42210 21375
rect 43710 21360 43890 21375
rect 5310 21225 5490 21240
rect 6990 21225 7170 21240
rect 5310 21210 7170 21225
rect 5310 21090 5340 21210
rect 5460 21090 7020 21210
rect 7140 21090 7170 21210
rect 5310 21075 7170 21090
rect 5310 21060 5490 21075
rect 6990 21060 7170 21075
rect 10110 21225 10290 21240
rect 11790 21225 11970 21240
rect 10110 21210 11970 21225
rect 10110 21090 10140 21210
rect 10260 21090 11820 21210
rect 11940 21090 11970 21210
rect 10110 21075 11970 21090
rect 10110 21060 10290 21075
rect 11790 21060 11970 21075
rect 17550 21225 17730 21240
rect 18270 21225 18450 21240
rect 17550 21210 18450 21225
rect 17550 21090 17580 21210
rect 17700 21090 18300 21210
rect 18420 21090 18450 21210
rect 17550 21075 18450 21090
rect 17550 21060 17730 21075
rect 18270 21060 18450 21075
rect 28830 21225 29010 21240
rect 29790 21225 29970 21240
rect 32670 21225 32850 21240
rect 28830 21210 32850 21225
rect 28830 21090 28860 21210
rect 28980 21090 29820 21210
rect 29940 21090 32700 21210
rect 32820 21090 32850 21210
rect 28830 21075 32850 21090
rect 28830 21060 29010 21075
rect 29790 21060 29970 21075
rect 32670 21060 32850 21075
rect 36750 21225 36930 21240
rect 42510 21225 42690 21240
rect 36750 21210 42690 21225
rect 36750 21090 36780 21210
rect 36900 21090 42540 21210
rect 42660 21090 42690 21210
rect 36750 21075 42690 21090
rect 44685 21225 44835 21375
rect 47310 21510 48210 21525
rect 47310 21390 47340 21510
rect 47460 21390 48060 21510
rect 48180 21390 48210 21510
rect 47310 21375 48210 21390
rect 47310 21360 47490 21375
rect 48030 21360 48210 21375
rect 45630 21225 45810 21240
rect 44685 21210 45810 21225
rect 44685 21090 45660 21210
rect 45780 21090 45810 21210
rect 44685 21075 45810 21090
rect 36750 21060 36930 21075
rect 42510 21060 42690 21075
rect 45630 21060 45810 21075
rect 6750 20925 6930 20940
rect 9630 20925 9810 20940
rect 6750 20910 9810 20925
rect 6750 20790 6780 20910
rect 6900 20790 9660 20910
rect 9780 20790 9810 20910
rect 6750 20775 9810 20790
rect 6750 20760 6930 20775
rect 9630 20760 9810 20775
rect 18510 20925 18690 20940
rect 20190 20925 20370 20940
rect 18510 20910 20370 20925
rect 18510 20790 18540 20910
rect 18660 20790 20220 20910
rect 20340 20790 20370 20910
rect 18510 20775 20370 20790
rect 18510 20760 18690 20775
rect 20190 20760 20370 20775
rect 40590 20925 40770 20940
rect 42270 20925 42450 20940
rect 42750 20925 42930 20940
rect 43710 20925 43890 20940
rect 40590 20910 43890 20925
rect 40590 20790 40620 20910
rect 40740 20790 42300 20910
rect 42420 20790 42780 20910
rect 42900 20790 43740 20910
rect 43860 20790 43890 20910
rect 40590 20775 43890 20790
rect 40590 20760 40770 20775
rect 42270 20760 42450 20775
rect 42750 20760 42930 20775
rect 43710 20760 43890 20775
rect 8910 20625 9090 20640
rect 11550 20625 11730 20640
rect 8910 20610 11730 20625
rect 8910 20490 8940 20610
rect 9060 20490 11580 20610
rect 11700 20490 11730 20610
rect 8910 20475 11730 20490
rect 8910 20460 9090 20475
rect 11550 20460 11730 20475
rect 19470 20625 19650 20640
rect 20430 20625 20610 20640
rect 19470 20610 20610 20625
rect 19470 20490 19500 20610
rect 19620 20490 20460 20610
rect 20580 20490 20610 20610
rect 19470 20475 20610 20490
rect 19470 20460 19650 20475
rect 20430 20460 20610 20475
rect 30510 20625 30690 20640
rect 31230 20625 31410 20640
rect 37470 20625 37650 20640
rect 30510 20610 37650 20625
rect 30510 20490 30540 20610
rect 30660 20490 31260 20610
rect 31380 20490 37500 20610
rect 37620 20490 37650 20610
rect 30510 20475 37650 20490
rect 30510 20460 30690 20475
rect 31230 20460 31410 20475
rect 37470 20460 37650 20475
rect 44910 20625 45090 20640
rect 49950 20625 50130 20640
rect 44910 20610 50130 20625
rect 44910 20490 44940 20610
rect 45060 20490 49980 20610
rect 50100 20490 50130 20610
rect 44910 20475 50130 20490
rect 44910 20460 45090 20475
rect 49950 20460 50130 20475
rect 15630 20325 15810 20340
rect 19710 20325 19890 20340
rect 15630 20310 19890 20325
rect 15630 20190 15660 20310
rect 15780 20190 19740 20310
rect 19860 20190 19890 20310
rect 15630 20175 19890 20190
rect 15630 20160 15810 20175
rect 19710 20160 19890 20175
rect 30990 20325 31170 20340
rect 45150 20325 45330 20340
rect 30990 20310 45330 20325
rect 30990 20190 31020 20310
rect 31140 20190 45180 20310
rect 45300 20190 45330 20310
rect 30990 20175 45330 20190
rect 30990 20160 31170 20175
rect 45150 20160 45330 20175
rect 24030 20025 24210 20040
rect 24510 20025 24690 20040
rect 24030 20010 24690 20025
rect 24030 19890 24060 20010
rect 24180 19890 24540 20010
rect 24660 19890 24690 20010
rect 24030 19875 24690 19890
rect 24030 19860 24210 19875
rect 24510 19860 24690 19875
rect 25950 20025 26130 20040
rect 30750 20025 30930 20040
rect 25950 20010 30930 20025
rect 25950 19890 25980 20010
rect 26100 19890 30780 20010
rect 30900 19890 30930 20010
rect 25950 19875 30930 19890
rect 25950 19860 26130 19875
rect 30750 19860 30930 19875
rect 36030 20025 36210 20040
rect 37470 20025 37650 20040
rect 36030 20010 37650 20025
rect 36030 19890 36060 20010
rect 36180 19890 37500 20010
rect 37620 19890 37650 20010
rect 36030 19875 37650 19890
rect 36030 19860 36210 19875
rect 37470 19860 37650 19875
rect 40350 20025 40530 20040
rect 42270 20025 42450 20040
rect 40350 20010 42450 20025
rect 40350 19890 40380 20010
rect 40500 19890 42300 20010
rect 42420 19890 42450 20010
rect 40350 19875 42450 19890
rect 40350 19860 40530 19875
rect 42270 19860 42450 19875
rect 46590 20025 46770 20040
rect 47550 20025 47730 20040
rect 46590 20010 47730 20025
rect 46590 19890 46620 20010
rect 46740 19890 47580 20010
rect 47700 19890 47730 20010
rect 46590 19875 47730 19890
rect 46590 19860 46770 19875
rect 47550 19860 47730 19875
rect 24510 19725 24690 19740
rect 26910 19725 27090 19740
rect 24510 19710 27090 19725
rect 24510 19590 24540 19710
rect 24660 19590 26940 19710
rect 27060 19590 27090 19710
rect 24510 19575 27090 19590
rect 24510 19560 24690 19575
rect 26910 19560 27090 19575
rect 33390 19725 33570 19740
rect 35070 19725 35250 19740
rect 33390 19710 35250 19725
rect 33390 19590 33420 19710
rect 33540 19590 35100 19710
rect 35220 19590 35250 19710
rect 33390 19575 35250 19590
rect 33390 19560 33570 19575
rect 35070 19560 35250 19575
rect 36510 19725 36690 19740
rect 37230 19725 37410 19740
rect 36510 19710 37410 19725
rect 36510 19590 36540 19710
rect 36660 19590 37260 19710
rect 37380 19590 37410 19710
rect 36510 19575 37410 19590
rect 36510 19560 36690 19575
rect 37230 19560 37410 19575
rect 41550 19725 41730 19740
rect 42030 19725 42210 19740
rect 41550 19710 42210 19725
rect 41550 19590 41580 19710
rect 41700 19590 42060 19710
rect 42180 19590 42210 19710
rect 41550 19575 42210 19590
rect 41550 19560 41730 19575
rect 42030 19560 42210 19575
rect 13230 19425 13410 19440
rect 14910 19425 15090 19440
rect 13230 19410 15090 19425
rect 13230 19290 13260 19410
rect 13380 19290 14940 19410
rect 15060 19290 15090 19410
rect 13230 19275 15090 19290
rect 13230 19260 13410 19275
rect 14910 19260 15090 19275
rect 26190 19425 26370 19440
rect 27150 19425 27330 19440
rect 26190 19410 27330 19425
rect 26190 19290 26220 19410
rect 26340 19290 27180 19410
rect 27300 19290 27330 19410
rect 26190 19275 27330 19290
rect 26190 19260 26370 19275
rect 27150 19260 27330 19275
rect 34590 19425 34770 19440
rect 36510 19425 36690 19440
rect 34590 19410 36690 19425
rect 34590 19290 34620 19410
rect 34740 19290 36540 19410
rect 36660 19290 36690 19410
rect 34590 19275 36690 19290
rect 34590 19260 34770 19275
rect 36510 19260 36690 19275
rect 39630 19425 39810 19440
rect 41070 19425 41250 19440
rect 39630 19410 41250 19425
rect 39630 19290 39660 19410
rect 39780 19290 41100 19410
rect 41220 19290 41250 19410
rect 39630 19275 41250 19290
rect 39630 19260 39810 19275
rect 41070 19260 41250 19275
rect 47550 19425 47730 19440
rect 48030 19425 48210 19440
rect 47550 19410 48210 19425
rect 47550 19290 47580 19410
rect 47700 19290 48060 19410
rect 48180 19290 48210 19410
rect 47550 19275 48210 19290
rect 47550 19260 47730 19275
rect 48030 19260 48210 19275
rect 15390 19125 15570 19140
rect 18510 19125 18690 19140
rect 15390 19110 18690 19125
rect 15390 18990 15420 19110
rect 15540 18990 18540 19110
rect 18660 18990 18690 19110
rect 15390 18975 18690 18990
rect 15390 18960 15570 18975
rect 18510 18960 18690 18975
rect 22110 19125 22290 19140
rect 22590 19125 22770 19140
rect 22110 19110 22770 19125
rect 22110 18990 22140 19110
rect 22260 18990 22620 19110
rect 22740 18990 22770 19110
rect 22110 18975 22770 18990
rect 22110 18960 22290 18975
rect 22590 18960 22770 18975
rect 24270 19125 24450 19140
rect 26190 19125 26370 19140
rect 24270 19110 26370 19125
rect 24270 18990 24300 19110
rect 24420 18990 26220 19110
rect 26340 18990 26370 19110
rect 24270 18975 26370 18990
rect 24270 18960 24450 18975
rect 26190 18960 26370 18975
rect 29550 19125 29730 19140
rect 30990 19125 31170 19140
rect 29550 19110 31170 19125
rect 29550 18990 29580 19110
rect 29700 18990 31020 19110
rect 31140 18990 31170 19110
rect 29550 18975 31170 18990
rect 29550 18960 29730 18975
rect 30990 18960 31170 18975
rect 31950 19125 32130 19140
rect 36030 19125 36210 19140
rect 31950 19110 36210 19125
rect 31950 18990 31980 19110
rect 32100 18990 36060 19110
rect 36180 18990 36210 19110
rect 31950 18975 36210 18990
rect 31950 18960 32130 18975
rect 36030 18960 36210 18975
rect 38910 19125 39090 19140
rect 39390 19125 39570 19140
rect 38910 19110 39570 19125
rect 38910 18990 38940 19110
rect 39060 18990 39420 19110
rect 39540 18990 39570 19110
rect 38910 18975 39570 18990
rect 38910 18960 39090 18975
rect 39390 18960 39570 18975
rect 41790 19125 41970 19140
rect 43470 19125 43650 19140
rect 41790 19110 43650 19125
rect 41790 18990 41820 19110
rect 41940 18990 43500 19110
rect 43620 18990 43650 19110
rect 41790 18975 43650 18990
rect 41790 18960 41970 18975
rect 43470 18960 43650 18975
rect 44670 19125 44850 19140
rect 45390 19125 45570 19140
rect 44670 19110 45570 19125
rect 44670 18990 44700 19110
rect 44820 18990 45420 19110
rect 45540 18990 45570 19110
rect 44670 18975 45570 18990
rect 44670 18960 44850 18975
rect 45390 18960 45570 18975
rect 13470 18825 13650 18840
rect 15630 18825 15810 18840
rect 18270 18825 18450 18840
rect 13470 18810 18450 18825
rect 13470 18690 13500 18810
rect 13620 18690 15660 18810
rect 15780 18690 18300 18810
rect 18420 18690 18450 18810
rect 13470 18675 18450 18690
rect 13470 18660 13650 18675
rect 15630 18660 15810 18675
rect 18270 18660 18450 18675
rect 20910 18825 21090 18840
rect 22830 18825 23010 18840
rect 20910 18810 23010 18825
rect 20910 18690 20940 18810
rect 21060 18690 22860 18810
rect 22980 18690 23010 18810
rect 20910 18675 23010 18690
rect 20910 18660 21090 18675
rect 22830 18660 23010 18675
rect 26430 18825 26610 18840
rect 26910 18825 27090 18840
rect 26430 18810 27090 18825
rect 26430 18690 26460 18810
rect 26580 18690 26940 18810
rect 27060 18690 27090 18810
rect 26430 18675 27090 18690
rect 26430 18660 26610 18675
rect 26910 18660 27090 18675
rect 31950 18825 32130 18840
rect 33630 18825 33810 18840
rect 31950 18810 33810 18825
rect 31950 18690 31980 18810
rect 32100 18690 33660 18810
rect 33780 18690 33810 18810
rect 31950 18675 33810 18690
rect 31950 18660 32130 18675
rect 33630 18660 33810 18675
rect 35550 18825 35730 18840
rect 43950 18825 44130 18840
rect 35550 18810 44130 18825
rect 35550 18690 35580 18810
rect 35700 18690 43980 18810
rect 44100 18690 44130 18810
rect 35550 18675 44130 18690
rect 35550 18660 35730 18675
rect 43950 18660 44130 18675
rect 44430 18825 44610 18840
rect 46590 18825 46770 18840
rect 44430 18810 46770 18825
rect 44430 18690 44460 18810
rect 44580 18690 46620 18810
rect 46740 18690 46770 18810
rect 44430 18675 46770 18690
rect 44430 18660 44610 18675
rect 46590 18660 46770 18675
rect 11550 18525 11730 18540
rect 17310 18525 17490 18540
rect 11550 18510 17490 18525
rect 11550 18390 11580 18510
rect 11700 18390 17340 18510
rect 17460 18390 17490 18510
rect 11550 18375 17490 18390
rect 11550 18360 11730 18375
rect 17310 18360 17490 18375
rect 20910 18525 21090 18540
rect 21390 18525 21570 18540
rect 20910 18510 21570 18525
rect 20910 18390 20940 18510
rect 21060 18390 21420 18510
rect 21540 18390 21570 18510
rect 20910 18375 21570 18390
rect 20910 18360 21090 18375
rect 21390 18360 21570 18375
rect 28350 18525 28530 18540
rect 29310 18525 29490 18540
rect 28350 18510 29490 18525
rect 28350 18390 28380 18510
rect 28500 18390 29340 18510
rect 29460 18390 29490 18510
rect 28350 18375 29490 18390
rect 28350 18360 28530 18375
rect 29310 18360 29490 18375
rect 32910 18525 33090 18540
rect 33630 18525 33810 18540
rect 32910 18510 33810 18525
rect 32910 18390 32940 18510
rect 33060 18390 33660 18510
rect 33780 18390 33810 18510
rect 32910 18375 33810 18390
rect 32910 18360 33090 18375
rect 33630 18360 33810 18375
rect 36750 18525 36930 18540
rect 38430 18525 38610 18540
rect 36750 18510 38610 18525
rect 36750 18390 36780 18510
rect 36900 18390 38460 18510
rect 38580 18390 38610 18510
rect 36750 18375 38610 18390
rect 36750 18360 36930 18375
rect 38430 18360 38610 18375
rect 40350 18525 40530 18540
rect 43230 18525 43410 18540
rect 40350 18510 43410 18525
rect 40350 18390 40380 18510
rect 40500 18390 43260 18510
rect 43380 18390 43410 18510
rect 40350 18375 43410 18390
rect 40350 18360 40530 18375
rect 43230 18360 43410 18375
rect 46590 18525 46770 18540
rect 49710 18525 49890 18540
rect 46590 18510 49890 18525
rect 46590 18390 46620 18510
rect 46740 18390 49740 18510
rect 49860 18390 49890 18510
rect 46590 18375 49890 18390
rect 46590 18360 46770 18375
rect 49710 18360 49890 18375
rect 27390 18225 27570 18240
rect 38910 18225 39090 18240
rect 25965 18210 39090 18225
rect 25965 18090 27420 18210
rect 27540 18090 38940 18210
rect 39060 18090 39090 18210
rect 25965 18075 39090 18090
rect 19470 17925 19650 17940
rect 25965 17925 26115 18075
rect 27390 18060 27570 18075
rect 38910 18060 39090 18075
rect 19470 17910 26115 17925
rect 19470 17790 19500 17910
rect 19620 17790 26115 17910
rect 19470 17775 26115 17790
rect 33630 17925 33810 17940
rect 40830 17925 41010 17940
rect 33630 17910 41010 17925
rect 33630 17790 33660 17910
rect 33780 17790 40860 17910
rect 40980 17790 41010 17910
rect 33630 17775 41010 17790
rect 19470 17760 19650 17775
rect 33630 17760 33810 17775
rect 40830 17760 41010 17775
rect 10830 17625 11010 17640
rect 16110 17625 16290 17640
rect 10830 17610 16290 17625
rect 10830 17490 10860 17610
rect 10980 17490 16140 17610
rect 16260 17490 16290 17610
rect 10830 17475 16290 17490
rect 10830 17460 11010 17475
rect 16110 17460 16290 17475
rect 18270 17625 18450 17640
rect 25230 17625 25410 17640
rect 18270 17610 25410 17625
rect 18270 17490 18300 17610
rect 18420 17490 25260 17610
rect 25380 17490 25410 17610
rect 18270 17475 25410 17490
rect 18270 17460 18450 17475
rect 25230 17460 25410 17475
rect 37230 17625 37410 17640
rect 46830 17625 47010 17640
rect 37230 17610 47010 17625
rect 37230 17490 37260 17610
rect 37380 17490 46860 17610
rect 46980 17490 47010 17610
rect 37230 17475 47010 17490
rect 37230 17460 37410 17475
rect 46830 17460 47010 17475
rect 23550 17025 23730 17040
rect 24270 17025 24450 17040
rect 27870 17025 28050 17040
rect 35790 17025 35970 17040
rect 23550 17010 35970 17025
rect 23550 16890 23580 17010
rect 23700 16890 24300 17010
rect 24420 16890 27900 17010
rect 28020 16890 35820 17010
rect 35940 16890 35970 17010
rect 23550 16875 35970 16890
rect 23550 16860 23730 16875
rect 24270 16860 24450 16875
rect 27870 16860 28050 16875
rect 35790 16860 35970 16875
rect 8430 16725 8610 16740
rect 6285 16710 8610 16725
rect 6285 16590 8460 16710
rect 8580 16590 8610 16710
rect 6285 16575 8610 16590
rect 0 16425 6435 16575
rect 8430 16560 8610 16575
rect 24030 16725 24210 16740
rect 24750 16725 24930 16740
rect 24030 16710 24930 16725
rect 24030 16590 24060 16710
rect 24180 16590 24780 16710
rect 24900 16590 24930 16710
rect 24030 16575 24930 16590
rect 24030 16560 24210 16575
rect 24750 16560 24930 16575
rect 25950 16725 26130 16740
rect 26430 16725 26610 16740
rect 25950 16710 26610 16725
rect 25950 16590 25980 16710
rect 26100 16590 26460 16710
rect 26580 16590 26610 16710
rect 25950 16575 26610 16590
rect 25950 16560 26130 16575
rect 26430 16560 26610 16575
rect 9390 16425 9570 16440
rect 13950 16425 14130 16440
rect 27630 16425 27810 16440
rect 28350 16425 28530 16440
rect 9390 16410 14130 16425
rect 9390 16290 9420 16410
rect 9540 16290 13980 16410
rect 14100 16290 14130 16410
rect 9390 16275 14130 16290
rect 9390 16260 9570 16275
rect 13950 16260 14130 16275
rect 24045 16410 28530 16425
rect 24045 16290 27660 16410
rect 27780 16290 28380 16410
rect 28500 16290 28530 16410
rect 24045 16275 28530 16290
rect 2430 16125 2610 16140
rect 12510 16125 12690 16140
rect 16350 16125 16530 16140
rect 2430 16110 16530 16125
rect 2430 15990 2460 16110
rect 2580 15990 12540 16110
rect 12660 15990 16380 16110
rect 16500 15990 16530 16110
rect 2430 15975 16530 15990
rect 2430 15960 2610 15975
rect 12510 15960 12690 15975
rect 16350 15960 16530 15975
rect 20430 16125 20610 16140
rect 24045 16125 24195 16275
rect 27630 16260 27810 16275
rect 28350 16260 28530 16275
rect 20430 16110 24195 16125
rect 20430 15990 20460 16110
rect 20580 15990 24195 16110
rect 20430 15975 24195 15990
rect 24510 16125 24690 16140
rect 25230 16125 25410 16140
rect 24510 16110 25410 16125
rect 24510 15990 24540 16110
rect 24660 15990 25260 16110
rect 25380 15990 25410 16110
rect 24510 15975 25410 15990
rect 20430 15960 20610 15975
rect 24510 15960 24690 15975
rect 25230 15960 25410 15975
rect 32910 16125 33090 16140
rect 37950 16125 38130 16140
rect 39390 16125 39570 16140
rect 32910 16110 39570 16125
rect 32910 15990 32940 16110
rect 33060 15990 37980 16110
rect 38100 15990 39420 16110
rect 39540 15990 39570 16110
rect 32910 15975 39570 15990
rect 32910 15960 33090 15975
rect 37950 15960 38130 15975
rect 39390 15960 39570 15975
rect 6750 15825 6930 15840
rect 9390 15825 9570 15840
rect 6750 15810 9570 15825
rect 6750 15690 6780 15810
rect 6900 15690 9420 15810
rect 9540 15690 9570 15810
rect 6750 15675 9570 15690
rect 6750 15660 6930 15675
rect 9390 15660 9570 15675
rect 12990 15825 13170 15840
rect 14190 15825 14370 15840
rect 12990 15810 14370 15825
rect 12990 15690 13020 15810
rect 13140 15690 14220 15810
rect 14340 15690 14370 15810
rect 12990 15675 14370 15690
rect 12990 15660 13170 15675
rect 14190 15660 14370 15675
rect 14910 15825 15090 15840
rect 16830 15825 17010 15840
rect 18510 15825 18690 15840
rect 21390 15825 21570 15840
rect 14910 15810 21570 15825
rect 14910 15690 14940 15810
rect 15060 15690 16860 15810
rect 16980 15690 18540 15810
rect 18660 15690 21420 15810
rect 21540 15690 21570 15810
rect 14910 15675 21570 15690
rect 14910 15660 15090 15675
rect 16830 15660 17010 15675
rect 18510 15660 18690 15675
rect 21390 15660 21570 15675
rect 22110 15825 22290 15840
rect 24990 15825 25170 15840
rect 22110 15810 25170 15825
rect 22110 15690 22140 15810
rect 22260 15690 25020 15810
rect 25140 15690 25170 15810
rect 22110 15675 25170 15690
rect 22110 15660 22290 15675
rect 24990 15660 25170 15675
rect 30030 15825 30210 15840
rect 31950 15825 32130 15840
rect 30030 15810 32130 15825
rect 30030 15690 30060 15810
rect 30180 15690 31980 15810
rect 32100 15690 32130 15810
rect 30030 15675 32130 15690
rect 30030 15660 30210 15675
rect 31950 15660 32130 15675
rect 35790 15825 35970 15840
rect 36270 15825 36450 15840
rect 35790 15810 36450 15825
rect 35790 15690 35820 15810
rect 35940 15690 36300 15810
rect 36420 15690 36450 15810
rect 35790 15675 36450 15690
rect 35790 15660 35970 15675
rect 36270 15660 36450 15675
rect 42270 15825 42450 15840
rect 43710 15825 43890 15840
rect 42270 15810 43890 15825
rect 42270 15690 42300 15810
rect 42420 15690 43740 15810
rect 43860 15690 43890 15810
rect 42270 15675 43890 15690
rect 42270 15660 42450 15675
rect 43710 15660 43890 15675
rect 44430 15825 44610 15840
rect 46590 15825 46770 15840
rect 44430 15810 46770 15825
rect 44430 15690 44460 15810
rect 44580 15690 46620 15810
rect 46740 15690 46770 15810
rect 44430 15675 46770 15690
rect 44430 15660 44610 15675
rect 46590 15660 46770 15675
rect 9150 15525 9330 15540
rect 10110 15525 10290 15540
rect 9150 15510 10290 15525
rect 9150 15390 9180 15510
rect 9300 15390 10140 15510
rect 10260 15390 10290 15510
rect 9150 15375 10290 15390
rect 9150 15360 9330 15375
rect 10110 15360 10290 15375
rect 14670 15525 14850 15540
rect 15630 15525 15810 15540
rect 14670 15510 15810 15525
rect 14670 15390 14700 15510
rect 14820 15390 15660 15510
rect 15780 15390 15810 15510
rect 14670 15375 15810 15390
rect 14670 15360 14850 15375
rect 15630 15360 15810 15375
rect 22590 15525 22770 15540
rect 24030 15525 24210 15540
rect 25470 15525 25650 15540
rect 22590 15510 25650 15525
rect 22590 15390 22620 15510
rect 22740 15390 24060 15510
rect 24180 15390 25500 15510
rect 25620 15390 25650 15510
rect 22590 15375 25650 15390
rect 22590 15360 22770 15375
rect 24030 15360 24210 15375
rect 25470 15360 25650 15375
rect 34590 15525 34770 15540
rect 35310 15525 35490 15540
rect 34590 15510 35490 15525
rect 34590 15390 34620 15510
rect 34740 15390 35340 15510
rect 35460 15390 35490 15510
rect 34590 15375 35490 15390
rect 34590 15360 34770 15375
rect 35310 15360 35490 15375
rect 36270 15525 36450 15540
rect 38190 15525 38370 15540
rect 36270 15510 38370 15525
rect 36270 15390 36300 15510
rect 36420 15390 38220 15510
rect 38340 15390 38370 15510
rect 36270 15375 38370 15390
rect 36270 15360 36450 15375
rect 38190 15360 38370 15375
rect 41310 15525 41490 15540
rect 42270 15525 42450 15540
rect 41310 15510 42450 15525
rect 41310 15390 41340 15510
rect 41460 15390 42300 15510
rect 42420 15390 42450 15510
rect 41310 15375 42450 15390
rect 41310 15360 41490 15375
rect 42270 15360 42450 15375
rect 49230 15525 49410 15540
rect 49710 15525 49890 15540
rect 49230 15510 49890 15525
rect 49230 15390 49260 15510
rect 49380 15390 49740 15510
rect 49860 15390 49890 15510
rect 49230 15375 49890 15390
rect 49230 15360 49410 15375
rect 49710 15360 49890 15375
rect 6030 15225 6210 15240
rect 10830 15225 11010 15240
rect 6030 15210 11010 15225
rect 6030 15090 6060 15210
rect 6180 15090 10860 15210
rect 10980 15090 11010 15210
rect 6030 15075 11010 15090
rect 6030 15060 6210 15075
rect 10830 15060 11010 15075
rect 16590 15225 16770 15240
rect 18750 15225 18930 15240
rect 20190 15225 20370 15240
rect 16590 15210 20370 15225
rect 16590 15090 16620 15210
rect 16740 15090 18780 15210
rect 18900 15090 20220 15210
rect 20340 15090 20370 15210
rect 16590 15075 20370 15090
rect 16590 15060 16770 15075
rect 18750 15060 18930 15075
rect 20190 15060 20370 15075
rect 23550 15225 23730 15240
rect 27150 15225 27330 15240
rect 23550 15210 27330 15225
rect 23550 15090 23580 15210
rect 23700 15090 27180 15210
rect 27300 15090 27330 15210
rect 23550 15075 27330 15090
rect 23550 15060 23730 15075
rect 27150 15060 27330 15075
rect 32430 15225 32610 15240
rect 35070 15225 35250 15240
rect 32430 15210 35250 15225
rect 32430 15090 32460 15210
rect 32580 15090 35100 15210
rect 35220 15090 35250 15210
rect 32430 15075 35250 15090
rect 32430 15060 32610 15075
rect 35070 15060 35250 15075
rect 36030 15225 36210 15240
rect 36990 15225 37170 15240
rect 36030 15210 37170 15225
rect 36030 15090 36060 15210
rect 36180 15090 37020 15210
rect 37140 15090 37170 15210
rect 36030 15075 37170 15090
rect 36030 15060 36210 15075
rect 36990 15060 37170 15075
rect 38190 15225 38370 15240
rect 42990 15225 43170 15240
rect 38190 15210 43170 15225
rect 38190 15090 38220 15210
rect 38340 15090 43020 15210
rect 43140 15090 43170 15210
rect 38190 15075 43170 15090
rect 38190 15060 38370 15075
rect 42990 15060 43170 15075
rect 44670 15225 44850 15240
rect 45390 15225 45570 15240
rect 49470 15225 49650 15240
rect 44670 15210 49650 15225
rect 44670 15090 44700 15210
rect 44820 15090 45420 15210
rect 45540 15090 49500 15210
rect 49620 15090 49650 15210
rect 44670 15075 49650 15090
rect 44670 15060 44850 15075
rect 45390 15060 45570 15075
rect 49470 15060 49650 15075
rect 11550 14925 11730 14940
rect 12510 14925 12690 14940
rect 11550 14910 12690 14925
rect 11550 14790 11580 14910
rect 11700 14790 12540 14910
rect 12660 14790 12690 14910
rect 11550 14775 12690 14790
rect 11550 14760 11730 14775
rect 12510 14760 12690 14775
rect 13710 14925 13890 14940
rect 17790 14925 17970 14940
rect 21870 14925 22050 14940
rect 13710 14910 22050 14925
rect 13710 14790 13740 14910
rect 13860 14790 17820 14910
rect 17940 14790 21900 14910
rect 22020 14790 22050 14910
rect 13710 14775 22050 14790
rect 13710 14760 13890 14775
rect 17790 14760 17970 14775
rect 21870 14760 22050 14775
rect 32670 14925 32850 14940
rect 33150 14925 33330 14940
rect 32670 14910 33330 14925
rect 32670 14790 32700 14910
rect 32820 14790 33180 14910
rect 33300 14790 33330 14910
rect 32670 14775 33330 14790
rect 32670 14760 32850 14775
rect 33150 14760 33330 14775
rect 35550 14925 35730 14940
rect 36270 14925 36450 14940
rect 35550 14910 36450 14925
rect 35550 14790 35580 14910
rect 35700 14790 36300 14910
rect 36420 14790 36450 14910
rect 35550 14775 36450 14790
rect 35550 14760 35730 14775
rect 36270 14760 36450 14775
rect 37710 14925 37890 14940
rect 41550 14925 41730 14940
rect 37710 14910 41730 14925
rect 37710 14790 37740 14910
rect 37860 14790 41580 14910
rect 41700 14790 41730 14910
rect 37710 14775 41730 14790
rect 37710 14760 37890 14775
rect 41550 14760 41730 14775
rect 43230 14925 43410 14940
rect 48030 14925 48210 14940
rect 43230 14910 48210 14925
rect 43230 14790 43260 14910
rect 43380 14790 48060 14910
rect 48180 14790 48210 14910
rect 43230 14775 48210 14790
rect 43230 14760 43410 14775
rect 48030 14760 48210 14775
rect 9630 14625 9810 14640
rect 11790 14625 11970 14640
rect 9630 14610 11970 14625
rect 9630 14490 9660 14610
rect 9780 14490 11820 14610
rect 11940 14490 11970 14610
rect 9630 14475 11970 14490
rect 9630 14460 9810 14475
rect 11790 14460 11970 14475
rect 16590 14625 16770 14640
rect 17070 14625 17250 14640
rect 16590 14610 17250 14625
rect 16590 14490 16620 14610
rect 16740 14490 17100 14610
rect 17220 14490 17250 14610
rect 16590 14475 17250 14490
rect 16590 14460 16770 14475
rect 17070 14460 17250 14475
rect 35790 14625 35970 14640
rect 39390 14625 39570 14640
rect 35790 14610 39570 14625
rect 35790 14490 35820 14610
rect 35940 14490 39420 14610
rect 39540 14490 39570 14610
rect 35790 14475 39570 14490
rect 35790 14460 35970 14475
rect 39390 14460 39570 14475
rect 11070 14325 11250 14340
rect 11550 14325 11730 14340
rect 11070 14310 11730 14325
rect 11070 14190 11100 14310
rect 11220 14190 11580 14310
rect 11700 14190 11730 14310
rect 11070 14175 11730 14190
rect 11070 14160 11250 14175
rect 11550 14160 11730 14175
rect 12750 14325 12930 14340
rect 19470 14325 19650 14340
rect 12750 14310 19650 14325
rect 12750 14190 12780 14310
rect 12900 14190 19500 14310
rect 19620 14190 19650 14310
rect 12750 14175 19650 14190
rect 12750 14160 12930 14175
rect 19470 14160 19650 14175
rect 34350 14325 34530 14340
rect 42510 14325 42690 14340
rect 34350 14310 42690 14325
rect 34350 14190 34380 14310
rect 34500 14190 42540 14310
rect 42660 14190 42690 14310
rect 34350 14175 42690 14190
rect 34350 14160 34530 14175
rect 42510 14160 42690 14175
rect 16830 14025 17010 14040
rect 17550 14025 17730 14040
rect 16830 14010 17730 14025
rect 16830 13890 16860 14010
rect 16980 13890 17580 14010
rect 17700 13890 17730 14010
rect 16830 13875 17730 13890
rect 16830 13860 17010 13875
rect 17550 13860 17730 13875
rect 31710 14025 31890 14040
rect 48270 14025 48450 14040
rect 31710 14010 48450 14025
rect 31710 13890 31740 14010
rect 31860 13890 48300 14010
rect 48420 13890 48450 14010
rect 31710 13875 48450 13890
rect 31710 13860 31890 13875
rect 48270 13860 48450 13875
rect 6990 13725 7170 13740
rect 18030 13725 18210 13740
rect 6990 13710 18210 13725
rect 6990 13590 7020 13710
rect 7140 13590 18060 13710
rect 18180 13590 18210 13710
rect 6990 13575 18210 13590
rect 6990 13560 7170 13575
rect 18030 13560 18210 13575
rect 20190 13725 20370 13740
rect 35310 13725 35490 13740
rect 20190 13710 35490 13725
rect 20190 13590 20220 13710
rect 20340 13590 35340 13710
rect 35460 13590 35490 13710
rect 20190 13575 35490 13590
rect 20190 13560 20370 13575
rect 35310 13560 35490 13575
rect 2670 13425 2850 13440
rect 9870 13425 10050 13440
rect 2670 13410 10050 13425
rect 2670 13290 2700 13410
rect 2820 13290 9900 13410
rect 10020 13290 10050 13410
rect 2670 13275 10050 13290
rect 2670 13260 2850 13275
rect 9870 13260 10050 13275
rect 15870 13425 16050 13440
rect 20190 13425 20370 13440
rect 15870 13410 20370 13425
rect 15870 13290 15900 13410
rect 16020 13290 20220 13410
rect 20340 13290 20370 13410
rect 15870 13275 20370 13290
rect 15870 13260 16050 13275
rect 20190 13260 20370 13275
rect 22350 13425 22530 13440
rect 26670 13425 26850 13440
rect 22350 13410 26850 13425
rect 22350 13290 22380 13410
rect 22500 13290 26700 13410
rect 26820 13290 26850 13410
rect 22350 13275 26850 13290
rect 22350 13260 22530 13275
rect 26670 13260 26850 13275
rect 31470 13425 31650 13440
rect 31950 13425 32130 13440
rect 31470 13410 32130 13425
rect 31470 13290 31500 13410
rect 31620 13290 31980 13410
rect 32100 13290 32130 13410
rect 31470 13275 32130 13290
rect 31470 13260 31650 13275
rect 31950 13260 32130 13275
rect 34590 13425 34770 13440
rect 36510 13425 36690 13440
rect 34590 13410 36690 13425
rect 34590 13290 34620 13410
rect 34740 13290 36540 13410
rect 36660 13290 36690 13410
rect 34590 13275 36690 13290
rect 34590 13260 34770 13275
rect 36510 13260 36690 13275
rect 8190 13125 8370 13140
rect 9390 13125 9570 13140
rect 8190 13110 9570 13125
rect 8190 12990 8220 13110
rect 8340 12990 9420 13110
rect 9540 12990 9570 13110
rect 8190 12975 9570 12990
rect 8190 12960 8370 12975
rect 9390 12960 9570 12975
rect 10830 13125 11010 13140
rect 12750 13125 12930 13140
rect 10830 13110 12930 13125
rect 10830 12990 10860 13110
rect 10980 12990 12780 13110
rect 12900 12990 12930 13110
rect 10830 12975 12930 12990
rect 10830 12960 11010 12975
rect 12750 12960 12930 12975
rect 17070 13125 17250 13140
rect 18990 13125 19170 13140
rect 17070 13110 19170 13125
rect 17070 12990 17100 13110
rect 17220 12990 19020 13110
rect 19140 12990 19170 13110
rect 17070 12975 19170 12990
rect 17070 12960 17250 12975
rect 18990 12960 19170 12975
rect 24750 13125 24930 13140
rect 26190 13125 26370 13140
rect 24750 13110 26370 13125
rect 24750 12990 24780 13110
rect 24900 12990 26220 13110
rect 26340 12990 26370 13110
rect 24750 12975 26370 12990
rect 24750 12960 24930 12975
rect 26190 12960 26370 12975
rect 26670 13125 26850 13140
rect 29550 13125 29730 13140
rect 26670 13110 29730 13125
rect 26670 12990 26700 13110
rect 26820 12990 29580 13110
rect 29700 12990 29730 13110
rect 26670 12975 29730 12990
rect 26670 12960 26850 12975
rect 29550 12960 29730 12975
rect 31950 13125 32130 13140
rect 32430 13125 32610 13140
rect 31950 13110 32610 13125
rect 31950 12990 31980 13110
rect 32100 12990 32460 13110
rect 32580 12990 32610 13110
rect 31950 12975 32610 12990
rect 31950 12960 32130 12975
rect 32430 12960 32610 12975
rect 32910 13125 33090 13140
rect 34590 13125 34770 13140
rect 32910 13110 34770 13125
rect 32910 12990 32940 13110
rect 33060 12990 34620 13110
rect 34740 12990 34770 13110
rect 32910 12975 34770 12990
rect 32910 12960 33090 12975
rect 34590 12960 34770 12975
rect 36030 13125 36210 13140
rect 36750 13125 36930 13140
rect 36030 13110 36930 13125
rect 36030 12990 36060 13110
rect 36180 12990 36780 13110
rect 36900 12990 36930 13110
rect 36030 12975 36930 12990
rect 36030 12960 36210 12975
rect 36750 12960 36930 12975
rect 39390 13125 39570 13140
rect 40830 13125 41010 13140
rect 39390 13110 41010 13125
rect 39390 12990 39420 13110
rect 39540 12990 40860 13110
rect 40980 12990 41010 13110
rect 39390 12975 41010 12990
rect 39390 12960 39570 12975
rect 40830 12960 41010 12975
rect 44430 13125 44610 13140
rect 45390 13125 45570 13140
rect 44430 13110 45570 13125
rect 44430 12990 44460 13110
rect 44580 12990 45420 13110
rect 45540 12990 45570 13110
rect 44430 12975 45570 12990
rect 44430 12960 44610 12975
rect 45390 12960 45570 12975
rect 18990 12825 19170 12840
rect 21630 12825 21810 12840
rect 18990 12810 21810 12825
rect 18990 12690 19020 12810
rect 19140 12690 21660 12810
rect 21780 12690 21810 12810
rect 18990 12675 21810 12690
rect 18990 12660 19170 12675
rect 21630 12660 21810 12675
rect 25230 12825 25410 12840
rect 26910 12825 27090 12840
rect 25230 12810 27090 12825
rect 25230 12690 25260 12810
rect 25380 12690 26940 12810
rect 27060 12690 27090 12810
rect 25230 12675 27090 12690
rect 25230 12660 25410 12675
rect 26910 12660 27090 12675
rect 29070 12825 29250 12840
rect 30750 12825 30930 12840
rect 29070 12810 30930 12825
rect 29070 12690 29100 12810
rect 29220 12690 30780 12810
rect 30900 12690 30930 12810
rect 29070 12675 30930 12690
rect 29070 12660 29250 12675
rect 30750 12660 30930 12675
rect 34830 12825 35010 12840
rect 37950 12825 38130 12840
rect 34830 12810 38130 12825
rect 34830 12690 34860 12810
rect 34980 12690 37980 12810
rect 38100 12690 38130 12810
rect 34830 12675 38130 12690
rect 34830 12660 35010 12675
rect 37950 12660 38130 12675
rect 38670 12825 38850 12840
rect 40590 12825 40770 12840
rect 38670 12810 40770 12825
rect 38670 12690 38700 12810
rect 38820 12690 40620 12810
rect 40740 12690 40770 12810
rect 38670 12675 40770 12690
rect 38670 12660 38850 12675
rect 40590 12660 40770 12675
rect 43230 12825 43410 12840
rect 43710 12825 43890 12840
rect 43230 12810 43890 12825
rect 43230 12690 43260 12810
rect 43380 12690 43740 12810
rect 43860 12690 43890 12810
rect 43230 12675 43890 12690
rect 43230 12660 43410 12675
rect 43710 12660 43890 12675
rect 44430 12825 44610 12840
rect 46590 12825 46770 12840
rect 44430 12810 46770 12825
rect 44430 12690 44460 12810
rect 44580 12690 46620 12810
rect 46740 12690 46770 12810
rect 44430 12675 46770 12690
rect 44430 12660 44610 12675
rect 46590 12660 46770 12675
rect 50190 12675 50370 12690
rect 55200 12675 55350 12690
rect 50190 12660 55350 12675
rect 50190 12540 50220 12660
rect 50340 12540 55350 12660
rect 11310 12525 11490 12540
rect 12510 12525 12690 12540
rect 15150 12525 15330 12540
rect 11310 12510 15330 12525
rect 11310 12390 11340 12510
rect 11460 12390 12540 12510
rect 12660 12390 15180 12510
rect 15300 12390 15330 12510
rect 11310 12375 15330 12390
rect 11310 12360 11490 12375
rect 12510 12360 12690 12375
rect 15150 12360 15330 12375
rect 21390 12525 21570 12540
rect 22590 12525 22770 12540
rect 21390 12510 22770 12525
rect 21390 12390 21420 12510
rect 21540 12390 22620 12510
rect 22740 12390 22770 12510
rect 21390 12375 22770 12390
rect 21390 12360 21570 12375
rect 22590 12360 22770 12375
rect 30270 12525 30450 12540
rect 32190 12525 32370 12540
rect 30270 12510 32370 12525
rect 30270 12390 30300 12510
rect 30420 12390 32220 12510
rect 32340 12390 32370 12510
rect 30270 12375 32370 12390
rect 30270 12360 30450 12375
rect 32190 12360 32370 12375
rect 37470 12525 37650 12540
rect 41070 12525 41250 12540
rect 37470 12510 41250 12525
rect 37470 12390 37500 12510
rect 37620 12390 41100 12510
rect 41220 12390 41250 12510
rect 37470 12375 41250 12390
rect 37470 12360 37650 12375
rect 41070 12360 41250 12375
rect 44670 12525 44850 12540
rect 46590 12525 46770 12540
rect 44670 12510 46770 12525
rect 44670 12390 44700 12510
rect 44820 12390 46620 12510
rect 46740 12390 46770 12510
rect 44670 12375 46770 12390
rect 44670 12360 44850 12375
rect 46590 12360 46770 12375
rect 47790 12525 47970 12540
rect 48270 12525 48450 12540
rect 48750 12525 48930 12540
rect 49230 12525 49410 12540
rect 47790 12510 49410 12525
rect 50190 12525 55350 12540
rect 50190 12510 50370 12525
rect 55200 12510 55350 12525
rect 47790 12390 47820 12510
rect 47940 12390 48300 12510
rect 48420 12390 48780 12510
rect 48900 12390 49260 12510
rect 49380 12390 49410 12510
rect 47790 12375 49410 12390
rect 47790 12360 47970 12375
rect 48270 12360 48450 12375
rect 48750 12360 48930 12375
rect 49230 12360 49410 12375
rect 30030 12225 30210 12240
rect 32190 12225 32370 12240
rect 30030 12210 32370 12225
rect 30030 12090 30060 12210
rect 30180 12090 32220 12210
rect 32340 12090 32370 12210
rect 30030 12075 32370 12090
rect 30030 12060 30210 12075
rect 32190 12060 32370 12075
rect 41550 12225 41730 12240
rect 48510 12225 48690 12240
rect 41550 12210 48690 12225
rect 41550 12090 41580 12210
rect 41700 12090 48540 12210
rect 48660 12090 48690 12210
rect 41550 12075 48690 12090
rect 41550 12060 41730 12075
rect 48510 12060 48690 12075
rect 24270 11925 24450 11940
rect 24750 11925 24930 11940
rect 24270 11910 24930 11925
rect 24270 11790 24300 11910
rect 24420 11790 24780 11910
rect 24900 11790 24930 11910
rect 24270 11775 24930 11790
rect 24270 11760 24450 11775
rect 24750 11760 24930 11775
rect 36270 11925 36450 11940
rect 43710 11925 43890 11940
rect 54510 11925 54690 11940
rect 36270 11910 54690 11925
rect 36270 11790 36300 11910
rect 36420 11790 43740 11910
rect 43860 11790 54540 11910
rect 54660 11790 54690 11910
rect 36270 11775 54690 11790
rect 36270 11760 36450 11775
rect 43710 11760 43890 11775
rect 54510 11760 54690 11775
rect 28350 11625 28530 11640
rect 50190 11625 50370 11640
rect 28350 11610 50370 11625
rect 28350 11490 28380 11610
rect 28500 11490 50220 11610
rect 50340 11490 50370 11610
rect 28350 11475 50370 11490
rect 28350 11460 28530 11475
rect 50190 11460 50370 11475
rect 5310 11175 5490 11190
rect 0 11160 5490 11175
rect 0 11040 5340 11160
rect 5460 11040 5490 11160
rect 0 11025 5490 11040
rect 5310 11010 5490 11025
rect 19950 11025 20130 11040
rect 20910 11025 21090 11040
rect 19950 11010 21090 11025
rect 19950 10890 19980 11010
rect 20100 10890 20940 11010
rect 21060 10890 21090 11010
rect 19950 10875 21090 10890
rect 19950 10860 20130 10875
rect 20910 10860 21090 10875
rect 15150 10725 15330 10740
rect 18030 10725 18210 10740
rect 15150 10710 18210 10725
rect 15150 10590 15180 10710
rect 15300 10590 18060 10710
rect 18180 10590 18210 10710
rect 15150 10575 18210 10590
rect 15150 10560 15330 10575
rect 18030 10560 18210 10575
rect 6270 10125 6450 10140
rect 7230 10125 7410 10140
rect 8430 10125 8610 10140
rect 6270 10110 8610 10125
rect 6270 9990 6300 10110
rect 6420 9990 7260 10110
rect 7380 9990 8460 10110
rect 8580 9990 8610 10110
rect 6270 9975 8610 9990
rect 6270 9960 6450 9975
rect 7230 9960 7410 9975
rect 8430 9960 8610 9975
rect 18750 10125 18930 10140
rect 19230 10125 19410 10140
rect 18750 10110 19410 10125
rect 18750 9990 18780 10110
rect 18900 9990 19260 10110
rect 19380 9990 19410 10110
rect 18750 9975 19410 9990
rect 18750 9960 18930 9975
rect 19230 9960 19410 9975
rect 31470 10125 31650 10140
rect 37230 10125 37410 10140
rect 41070 10125 41250 10140
rect 31470 10110 41250 10125
rect 31470 9990 31500 10110
rect 31620 9990 37260 10110
rect 37380 9990 41100 10110
rect 41220 9990 41250 10110
rect 31470 9975 41250 9990
rect 31470 9960 31650 9975
rect 37230 9960 37410 9975
rect 41070 9960 41250 9975
rect 5550 9825 5730 9840
rect 6510 9825 6690 9840
rect 5550 9810 6690 9825
rect 5550 9690 5580 9810
rect 5700 9690 6540 9810
rect 6660 9690 6690 9810
rect 5550 9675 6690 9690
rect 5550 9660 5730 9675
rect 6510 9660 6690 9675
rect 12510 9825 12690 9840
rect 23310 9825 23490 9840
rect 25470 9825 25650 9840
rect 12510 9810 25650 9825
rect 12510 9690 12540 9810
rect 12660 9690 23340 9810
rect 23460 9690 25500 9810
rect 25620 9690 25650 9810
rect 12510 9675 25650 9690
rect 12510 9660 12690 9675
rect 23310 9660 23490 9675
rect 25470 9660 25650 9675
rect 33150 9825 33330 9840
rect 33630 9825 33810 9840
rect 33150 9810 33810 9825
rect 33150 9690 33180 9810
rect 33300 9690 33660 9810
rect 33780 9690 33810 9810
rect 33150 9675 33810 9690
rect 33150 9660 33330 9675
rect 33630 9660 33810 9675
rect 36750 9825 36930 9840
rect 37470 9825 37650 9840
rect 38190 9825 38370 9840
rect 36750 9810 38370 9825
rect 36750 9690 36780 9810
rect 36900 9690 37500 9810
rect 37620 9690 38220 9810
rect 38340 9690 38370 9810
rect 36750 9675 38370 9690
rect 36750 9660 36930 9675
rect 37470 9660 37650 9675
rect 38190 9660 38370 9675
rect 42030 9825 42210 9840
rect 46830 9825 47010 9840
rect 42030 9810 47010 9825
rect 42030 9690 42060 9810
rect 42180 9690 46860 9810
rect 46980 9690 47010 9810
rect 42030 9675 47010 9690
rect 42030 9660 42210 9675
rect 46830 9660 47010 9675
rect 6750 9525 6930 9540
rect 8430 9525 8610 9540
rect 6750 9510 8610 9525
rect 6750 9390 6780 9510
rect 6900 9390 8460 9510
rect 8580 9390 8610 9510
rect 6750 9375 8610 9390
rect 6750 9360 6930 9375
rect 8430 9360 8610 9375
rect 9390 9525 9570 9540
rect 9870 9525 10050 9540
rect 10350 9525 10530 9540
rect 9390 9510 10530 9525
rect 9390 9390 9420 9510
rect 9540 9390 9900 9510
rect 10020 9390 10380 9510
rect 10500 9390 10530 9510
rect 9390 9375 10530 9390
rect 9390 9360 9570 9375
rect 9870 9360 10050 9375
rect 10350 9360 10530 9375
rect 16350 9525 16530 9540
rect 21870 9525 22050 9540
rect 16350 9510 22050 9525
rect 16350 9390 16380 9510
rect 16500 9390 21900 9510
rect 22020 9390 22050 9510
rect 16350 9375 22050 9390
rect 16350 9360 16530 9375
rect 21870 9360 22050 9375
rect 39150 9525 39330 9540
rect 39870 9525 40050 9540
rect 39150 9510 40050 9525
rect 39150 9390 39180 9510
rect 39300 9390 39900 9510
rect 40020 9390 40050 9510
rect 39150 9375 40050 9390
rect 39150 9360 39330 9375
rect 39870 9360 40050 9375
rect 7710 9225 7890 9240
rect 9630 9225 9810 9240
rect 10110 9225 10290 9240
rect 7710 9210 10290 9225
rect 7710 9090 7740 9210
rect 7860 9090 9660 9210
rect 9780 9090 10140 9210
rect 10260 9090 10290 9210
rect 7710 9075 10290 9090
rect 7710 9060 7890 9075
rect 9630 9060 9810 9075
rect 10110 9060 10290 9075
rect 16350 9225 16530 9240
rect 17310 9225 17490 9240
rect 16350 9210 17490 9225
rect 16350 9090 16380 9210
rect 16500 9090 17340 9210
rect 17460 9090 17490 9210
rect 16350 9075 17490 9090
rect 16350 9060 16530 9075
rect 17310 9060 17490 9075
rect 19230 9225 19410 9240
rect 20910 9225 21090 9240
rect 19230 9210 21090 9225
rect 19230 9090 19260 9210
rect 19380 9090 20940 9210
rect 21060 9090 21090 9210
rect 19230 9075 21090 9090
rect 19230 9060 19410 9075
rect 20910 9060 21090 9075
rect 21630 9225 21810 9240
rect 24030 9225 24210 9240
rect 21630 9210 24210 9225
rect 21630 9090 21660 9210
rect 21780 9090 24060 9210
rect 24180 9090 24210 9210
rect 21630 9075 24210 9090
rect 21630 9060 21810 9075
rect 24030 9060 24210 9075
rect 29550 9225 29730 9240
rect 30990 9225 31170 9240
rect 29550 9210 31170 9225
rect 29550 9090 29580 9210
rect 29700 9090 31020 9210
rect 31140 9090 31170 9210
rect 29550 9075 31170 9090
rect 29550 9060 29730 9075
rect 30990 9060 31170 9075
rect 32430 9225 32610 9240
rect 39390 9225 39570 9240
rect 32430 9210 39570 9225
rect 32430 9090 32460 9210
rect 32580 9090 39420 9210
rect 39540 9090 39570 9210
rect 32430 9075 39570 9090
rect 32430 9060 32610 9075
rect 39390 9060 39570 9075
rect 42270 9225 42450 9240
rect 43950 9225 44130 9240
rect 42270 9210 44130 9225
rect 42270 9090 42300 9210
rect 42420 9090 43980 9210
rect 44100 9090 44130 9210
rect 42270 9075 44130 9090
rect 42270 9060 42450 9075
rect 43950 9060 44130 9075
rect 47550 9225 47730 9240
rect 49470 9225 49650 9240
rect 47550 9210 49650 9225
rect 47550 9090 47580 9210
rect 47700 9090 49500 9210
rect 49620 9090 49650 9210
rect 47550 9075 49650 9090
rect 47550 9060 47730 9075
rect 49470 9060 49650 9075
rect 18990 8925 19170 8940
rect 20910 8925 21090 8940
rect 18990 8910 21090 8925
rect 18990 8790 19020 8910
rect 19140 8790 20940 8910
rect 21060 8790 21090 8910
rect 18990 8775 21090 8790
rect 18990 8760 19170 8775
rect 20910 8760 21090 8775
rect 23790 8925 23970 8940
rect 24510 8925 24690 8940
rect 28350 8925 28530 8940
rect 23790 8910 28530 8925
rect 23790 8790 23820 8910
rect 23940 8790 24540 8910
rect 24660 8790 28380 8910
rect 28500 8790 28530 8910
rect 23790 8775 28530 8790
rect 23790 8760 23970 8775
rect 24510 8760 24690 8775
rect 28350 8760 28530 8775
rect 29070 8925 29250 8940
rect 29790 8925 29970 8940
rect 29070 8910 29970 8925
rect 29070 8790 29100 8910
rect 29220 8790 29820 8910
rect 29940 8790 29970 8910
rect 29070 8775 29970 8790
rect 29070 8760 29250 8775
rect 29790 8760 29970 8775
rect 18750 8625 18930 8640
rect 21150 8625 21330 8640
rect 18750 8610 21330 8625
rect 18750 8490 18780 8610
rect 18900 8490 21180 8610
rect 21300 8490 21330 8610
rect 18750 8475 21330 8490
rect 18750 8460 18930 8475
rect 21150 8460 21330 8475
rect 28830 8625 29010 8640
rect 29550 8625 29730 8640
rect 28830 8610 29730 8625
rect 28830 8490 28860 8610
rect 28980 8490 29580 8610
rect 29700 8490 29730 8610
rect 28830 8475 29730 8490
rect 28830 8460 29010 8475
rect 29550 8460 29730 8475
rect 42510 8025 42690 8040
rect 48030 8025 48210 8040
rect 42510 8010 48210 8025
rect 42510 7890 42540 8010
rect 42660 7890 48060 8010
rect 48180 7890 48210 8010
rect 42510 7875 48210 7890
rect 42510 7860 42690 7875
rect 48030 7860 48210 7875
rect 17790 7725 17970 7740
rect 18510 7725 18690 7740
rect 17790 7710 18690 7725
rect 17790 7590 17820 7710
rect 17940 7590 18540 7710
rect 18660 7590 18690 7710
rect 17790 7575 18690 7590
rect 17790 7560 17970 7575
rect 18510 7560 18690 7575
rect 26430 7725 26610 7740
rect 26910 7725 27090 7740
rect 26430 7710 27090 7725
rect 26430 7590 26460 7710
rect 26580 7590 26940 7710
rect 27060 7590 27090 7710
rect 26430 7575 27090 7590
rect 26430 7560 26610 7575
rect 26910 7560 27090 7575
rect 28350 7725 28530 7740
rect 32670 7725 32850 7740
rect 35310 7725 35490 7740
rect 28350 7710 35490 7725
rect 28350 7590 28380 7710
rect 28500 7590 32700 7710
rect 32820 7590 35340 7710
rect 35460 7590 35490 7710
rect 28350 7575 35490 7590
rect 28350 7560 28530 7575
rect 32670 7560 32850 7575
rect 35310 7560 35490 7575
rect 36510 7725 36690 7740
rect 38430 7725 38610 7740
rect 40350 7725 40530 7740
rect 36510 7710 40530 7725
rect 36510 7590 36540 7710
rect 36660 7590 38460 7710
rect 38580 7590 40380 7710
rect 40500 7590 40530 7710
rect 36510 7575 40530 7590
rect 36510 7560 36690 7575
rect 38430 7560 38610 7575
rect 40350 7560 40530 7575
rect 40830 7725 41010 7740
rect 44910 7725 45090 7740
rect 40830 7710 45090 7725
rect 40830 7590 40860 7710
rect 40980 7590 44940 7710
rect 45060 7590 45090 7710
rect 40830 7575 45090 7590
rect 40830 7560 41010 7575
rect 44910 7560 45090 7575
rect 8190 7425 8370 7440
rect 10110 7425 10290 7440
rect 8190 7410 10290 7425
rect 8190 7290 8220 7410
rect 8340 7290 10140 7410
rect 10260 7290 10290 7410
rect 8190 7275 10290 7290
rect 8190 7260 8370 7275
rect 10110 7260 10290 7275
rect 26190 7425 26370 7440
rect 35070 7425 35250 7440
rect 36750 7425 36930 7440
rect 26190 7410 36930 7425
rect 26190 7290 26220 7410
rect 26340 7290 35100 7410
rect 35220 7290 36780 7410
rect 36900 7290 36930 7410
rect 26190 7275 36930 7290
rect 26190 7260 26370 7275
rect 35070 7260 35250 7275
rect 36750 7260 36930 7275
rect 37230 7425 37410 7440
rect 46590 7425 46770 7440
rect 47310 7425 47490 7440
rect 37230 7410 47490 7425
rect 37230 7290 37260 7410
rect 37380 7290 46620 7410
rect 46740 7290 47340 7410
rect 47460 7290 47490 7410
rect 37230 7275 47490 7290
rect 37230 7260 37410 7275
rect 46590 7260 46770 7275
rect 47310 7260 47490 7275
rect 5550 7125 5730 7140
rect 10350 7125 10530 7140
rect 5550 7110 10530 7125
rect 5550 6990 5580 7110
rect 5700 6990 10380 7110
rect 10500 6990 10530 7110
rect 5550 6975 10530 6990
rect 5550 6960 5730 6975
rect 10350 6960 10530 6975
rect 12270 7125 12450 7140
rect 12750 7125 12930 7140
rect 15870 7125 16050 7140
rect 12270 7110 16050 7125
rect 12270 6990 12300 7110
rect 12420 6990 12780 7110
rect 12900 6990 15900 7110
rect 16020 6990 16050 7110
rect 12270 6975 16050 6990
rect 12270 6960 12450 6975
rect 12750 6960 12930 6975
rect 15870 6960 16050 6975
rect 24270 7125 24450 7140
rect 27870 7125 28050 7140
rect 24270 7110 28050 7125
rect 24270 6990 24300 7110
rect 24420 6990 27900 7110
rect 28020 6990 28050 7110
rect 24270 6975 28050 6990
rect 24270 6960 24450 6975
rect 27870 6960 28050 6975
rect 30030 7125 30210 7140
rect 31710 7125 31890 7140
rect 32910 7125 33090 7140
rect 30030 7110 33090 7125
rect 30030 6990 30060 7110
rect 30180 6990 31740 7110
rect 31860 6990 32940 7110
rect 33060 6990 33090 7110
rect 30030 6975 33090 6990
rect 30030 6960 30210 6975
rect 31710 6960 31890 6975
rect 32910 6960 33090 6975
rect 38430 7125 38610 7140
rect 38910 7125 39090 7140
rect 40830 7125 41010 7140
rect 38430 7110 41010 7125
rect 38430 6990 38460 7110
rect 38580 6990 38940 7110
rect 39060 6990 40860 7110
rect 40980 6990 41010 7110
rect 38430 6975 41010 6990
rect 38430 6960 38610 6975
rect 38910 6960 39090 6975
rect 40830 6960 41010 6975
rect 44670 7125 44850 7140
rect 46590 7125 46770 7140
rect 44670 7110 46770 7125
rect 44670 6990 44700 7110
rect 44820 6990 46620 7110
rect 46740 6990 46770 7110
rect 44670 6975 46770 6990
rect 44670 6960 44850 6975
rect 46590 6960 46770 6975
rect 9870 6825 10050 6840
rect 14190 6825 14370 6840
rect 9870 6810 14370 6825
rect 9870 6690 9900 6810
rect 10020 6690 14220 6810
rect 14340 6690 14370 6810
rect 9870 6675 14370 6690
rect 9870 6660 10050 6675
rect 14190 6660 14370 6675
rect 27630 6825 27810 6840
rect 30750 6825 30930 6840
rect 27630 6810 30930 6825
rect 27630 6690 27660 6810
rect 27780 6690 30780 6810
rect 30900 6690 30930 6810
rect 27630 6675 30930 6690
rect 27630 6660 27810 6675
rect 30750 6660 30930 6675
rect 32190 6825 32370 6840
rect 33630 6825 33810 6840
rect 32190 6810 33810 6825
rect 32190 6690 32220 6810
rect 32340 6690 33660 6810
rect 33780 6690 33810 6810
rect 32190 6675 33810 6690
rect 32190 6660 32370 6675
rect 33630 6660 33810 6675
rect 38910 6825 39090 6840
rect 39390 6825 39570 6840
rect 38910 6810 39570 6825
rect 38910 6690 38940 6810
rect 39060 6690 39420 6810
rect 39540 6690 39570 6810
rect 38910 6675 39570 6690
rect 38910 6660 39090 6675
rect 39390 6660 39570 6675
rect 44190 6825 44370 6840
rect 45390 6825 45570 6840
rect 46830 6825 47010 6840
rect 44190 6810 47010 6825
rect 44190 6690 44220 6810
rect 44340 6690 45420 6810
rect 45540 6690 46860 6810
rect 46980 6690 47010 6810
rect 44190 6675 47010 6690
rect 44190 6660 44370 6675
rect 45390 6660 45570 6675
rect 46830 6660 47010 6675
rect 2670 6525 2850 6540
rect 9390 6525 9570 6540
rect 10350 6525 10530 6540
rect 2670 6510 10530 6525
rect 2670 6390 2700 6510
rect 2820 6390 9420 6510
rect 9540 6390 10380 6510
rect 10500 6390 10530 6510
rect 2670 6375 10530 6390
rect 2670 6360 2850 6375
rect 9390 6360 9570 6375
rect 10350 6360 10530 6375
rect 10830 6525 11010 6540
rect 11790 6525 11970 6540
rect 10830 6510 11970 6525
rect 10830 6390 10860 6510
rect 10980 6390 11820 6510
rect 11940 6390 11970 6510
rect 10830 6375 11970 6390
rect 10830 6360 11010 6375
rect 11790 6360 11970 6375
rect 12270 6525 12450 6540
rect 12750 6525 12930 6540
rect 13230 6525 13410 6540
rect 15390 6525 15570 6540
rect 12270 6510 15570 6525
rect 12270 6390 12300 6510
rect 12420 6390 12780 6510
rect 12900 6390 13260 6510
rect 13380 6390 15420 6510
rect 15540 6390 15570 6510
rect 12270 6375 15570 6390
rect 12270 6360 12450 6375
rect 12750 6360 12930 6375
rect 13230 6360 13410 6375
rect 15390 6360 15570 6375
rect 27870 6525 28050 6540
rect 28350 6525 28530 6540
rect 27870 6510 28530 6525
rect 27870 6390 27900 6510
rect 28020 6390 28380 6510
rect 28500 6390 28530 6510
rect 27870 6375 28530 6390
rect 27870 6360 28050 6375
rect 28350 6360 28530 6375
rect 30510 6525 30690 6540
rect 31470 6525 31650 6540
rect 30510 6510 31650 6525
rect 30510 6390 30540 6510
rect 30660 6390 31500 6510
rect 31620 6390 31650 6510
rect 30510 6375 31650 6390
rect 30510 6360 30690 6375
rect 31470 6360 31650 6375
rect 33150 6525 33330 6540
rect 34830 6525 35010 6540
rect 33150 6510 35010 6525
rect 33150 6390 33180 6510
rect 33300 6390 34860 6510
rect 34980 6390 35010 6510
rect 33150 6375 35010 6390
rect 33150 6360 33330 6375
rect 34830 6360 35010 6375
rect 37470 6525 37650 6540
rect 38430 6525 38610 6540
rect 37470 6510 38610 6525
rect 37470 6390 37500 6510
rect 37620 6390 38460 6510
rect 38580 6390 38610 6510
rect 37470 6375 38610 6390
rect 37470 6360 37650 6375
rect 38430 6360 38610 6375
rect 43950 6525 44130 6540
rect 47790 6525 47970 6540
rect 43950 6510 47970 6525
rect 43950 6390 43980 6510
rect 44100 6390 47820 6510
rect 47940 6390 47970 6510
rect 43950 6375 47970 6390
rect 43950 6360 44130 6375
rect 47790 6360 47970 6375
rect 6510 6225 6690 6240
rect 6990 6225 7170 6240
rect 6510 6210 7170 6225
rect 6510 6090 6540 6210
rect 6660 6090 7020 6210
rect 7140 6090 7170 6210
rect 6510 6075 7170 6090
rect 6510 6060 6690 6075
rect 6990 6060 7170 6075
rect 7710 6225 7890 6240
rect 12990 6225 13170 6240
rect 18510 6225 18690 6240
rect 7710 6210 18690 6225
rect 7710 6090 7740 6210
rect 7860 6090 13020 6210
rect 13140 6090 18540 6210
rect 18660 6090 18690 6210
rect 7710 6075 18690 6090
rect 7710 6060 7890 6075
rect 12990 6060 13170 6075
rect 18510 6060 18690 6075
rect 20670 6225 20850 6240
rect 32430 6225 32610 6240
rect 20670 6210 32610 6225
rect 20670 6090 20700 6210
rect 20820 6090 32460 6210
rect 32580 6090 32610 6210
rect 20670 6075 32610 6090
rect 20670 6060 20850 6075
rect 32430 6060 32610 6075
rect 36510 6225 36690 6240
rect 36990 6225 37170 6240
rect 36510 6210 37170 6225
rect 36510 6090 36540 6210
rect 36660 6090 37020 6210
rect 37140 6090 37170 6210
rect 36510 6075 37170 6090
rect 36510 6060 36690 6075
rect 36990 6060 37170 6075
rect 23310 5925 23490 5940
rect 27390 5925 27570 5940
rect 23310 5910 27570 5925
rect 23310 5790 23340 5910
rect 23460 5790 27420 5910
rect 27540 5790 27570 5910
rect 8430 5775 8610 5790
rect 0 5760 8610 5775
rect 23310 5775 27570 5790
rect 23310 5760 23490 5775
rect 27390 5760 27570 5775
rect 0 5640 8460 5760
rect 8580 5640 8610 5760
rect 0 5625 8610 5640
rect 8430 5610 8610 5625
rect 18510 5325 18690 5340
rect 50910 5325 51090 5340
rect 18510 5310 51090 5325
rect 18510 5190 18540 5310
rect 18660 5190 50940 5310
rect 51060 5190 51090 5310
rect 18510 5175 51090 5190
rect 18510 5160 18690 5175
rect 50910 5160 51090 5175
rect 54510 1155 54690 1170
rect 55200 1155 55350 1170
rect 54510 1140 55350 1155
rect 54510 1020 54540 1140
rect 54660 1020 55350 1140
rect 54510 1005 55350 1020
rect 54510 990 54690 1005
rect 55200 990 55350 1005
rect 12510 885 12690 900
rect 24750 885 24930 900
rect 12510 870 24930 885
rect 6270 855 6450 870
rect 0 840 6450 855
rect 0 720 6300 840
rect 6420 720 6450 840
rect 12510 750 12540 870
rect 12660 750 24780 870
rect 24900 750 24930 870
rect 12510 735 24930 750
rect 12510 720 12690 735
rect 24750 720 24930 735
rect 0 705 6450 720
rect 6270 690 6450 705
<< m1p >>
rect 11340 43290 11460 43410
rect 12780 43290 12900 43410
rect 21180 43290 21300 43410
rect 34620 43290 34740 43410
rect 41820 43290 41940 43410
rect 45420 43290 45540 43410
rect 5580 42990 5700 43110
rect 6300 42990 6420 43110
rect 6780 42990 6900 43110
rect 7740 42990 7860 43110
rect 8460 42990 8580 43110
rect 8940 42990 9060 43110
rect 10380 42990 10500 43110
rect 11100 42990 11220 43110
rect 12540 42990 12660 43110
rect 13740 42990 13860 43110
rect 14460 42990 14580 43110
rect 15420 42990 15540 43110
rect 17100 42990 17220 43110
rect 17820 42990 17940 43110
rect 19260 42990 19380 43110
rect 20700 42990 20820 43110
rect 21420 42990 21540 43110
rect 22620 42990 22740 43110
rect 24060 42990 24180 43110
rect 25020 42990 25140 43110
rect 25740 42990 25860 43110
rect 26700 42990 26820 43110
rect 27900 42990 28020 43110
rect 28620 42990 28740 43110
rect 29100 42990 29220 43110
rect 30300 42990 30420 43110
rect 31020 42990 31140 43110
rect 31740 42990 31860 43110
rect 32460 42990 32580 43110
rect 33660 42990 33780 43110
rect 34860 42990 34980 43110
rect 35820 42990 35940 43110
rect 37260 42990 37380 43110
rect 37740 42990 37860 43110
rect 38460 42990 38580 43110
rect 39420 42990 39540 43110
rect 40860 42990 40980 43110
rect 42060 42990 42180 43110
rect 43020 42990 43140 43110
rect 43740 42990 43860 43110
rect 44220 42990 44340 43110
rect 44940 42990 45060 43110
rect 45180 42990 45300 43110
rect 45660 42990 45780 43110
rect 47100 42990 47220 43110
rect 47340 42990 47460 43110
rect 48780 42990 48900 43110
rect 6060 42690 6180 42810
rect 7020 42690 7140 42810
rect 8220 42690 8340 42810
rect 9660 42690 9780 42810
rect 10860 42690 10980 42810
rect 12300 42690 12420 42810
rect 13980 42690 14100 42810
rect 15660 42690 15780 42810
rect 17340 42690 17460 42810
rect 19740 42690 19860 42810
rect 23340 42690 23460 42810
rect 25500 42690 25620 42810
rect 26940 42690 27060 42810
rect 28140 42690 28260 42810
rect 29340 42690 29460 42810
rect 30540 42690 30660 42810
rect 31980 42690 32100 42810
rect 33420 42690 33540 42810
rect 35100 42690 35220 42810
rect 36540 42690 36660 42810
rect 38220 42690 38340 42810
rect 40140 42690 40260 42810
rect 43260 42690 43380 42810
rect 44460 42690 44580 42810
rect 46380 42690 46500 42810
rect 48060 42690 48180 42810
rect 5580 42390 5700 42510
rect 7260 42390 7380 42510
rect 7740 42390 7860 42510
rect 14460 42390 14580 42510
rect 15900 42390 16020 42510
rect 17820 42390 17940 42510
rect 25020 42390 25140 42510
rect 27180 42390 27300 42510
rect 28620 42390 28740 42510
rect 29580 42390 29700 42510
rect 31020 42390 31140 42510
rect 32460 42390 32580 42510
rect 33180 42390 33300 42510
rect 37740 42390 37860 42510
rect 43740 42390 43860 42510
rect 44940 42390 45060 42510
rect 14460 39990 14580 40110
rect 8220 39690 8340 39810
rect 10140 39690 10260 39810
rect 13980 39690 14100 39810
rect 14940 39690 15060 39810
rect 17100 39690 17220 39810
rect 17580 39690 17700 39810
rect 19980 39690 20100 39810
rect 20940 39690 21060 39810
rect 25500 39690 25620 39810
rect 30540 39690 30660 39810
rect 31980 39690 32100 39810
rect 36780 39690 36900 39810
rect 37740 39690 37860 39810
rect 39660 39690 39780 39810
rect 40860 39690 40980 39810
rect 43740 39690 43860 39810
rect 45900 39690 46020 39810
rect 48300 39690 48420 39810
rect 49260 39690 49380 39810
rect 5820 39390 5940 39510
rect 6540 39390 6660 39510
rect 8460 39390 8580 39510
rect 9900 39390 10020 39510
rect 10620 39390 10740 39510
rect 11340 39390 11460 39510
rect 12540 39390 12660 39510
rect 13740 39390 13860 39510
rect 16620 39390 16740 39510
rect 18060 39390 18180 39510
rect 19500 39390 19620 39510
rect 21180 39390 21300 39510
rect 22620 39390 22740 39510
rect 24300 39390 24420 39510
rect 25020 39390 25140 39510
rect 26220 39390 26340 39510
rect 26700 39390 26820 39510
rect 27180 39390 27300 39510
rect 30780 39390 30900 39510
rect 32220 39390 32340 39510
rect 34140 39390 34260 39510
rect 36300 39390 36420 39510
rect 37980 39390 38100 39510
rect 39180 39390 39300 39510
rect 40620 39390 40740 39510
rect 43260 39390 43380 39510
rect 46380 39390 46500 39510
rect 47820 39390 47940 39510
rect 49500 39390 49620 39510
rect 6060 39090 6180 39210
rect 8700 39090 8820 39210
rect 9660 39090 9780 39210
rect 11100 39090 11220 39210
rect 11580 39090 11700 39210
rect 13020 39090 13140 39210
rect 13500 39090 13620 39210
rect 15180 39090 15300 39210
rect 15900 39090 16020 39210
rect 16380 39090 16500 39210
rect 17100 39090 17220 39210
rect 17580 39090 17700 39210
rect 18300 39090 18420 39210
rect 18540 39090 18660 39210
rect 19260 39090 19380 39210
rect 19980 39090 20100 39210
rect 21420 39090 21540 39210
rect 21900 39090 22020 39210
rect 23340 39090 23460 39210
rect 24060 39090 24180 39210
rect 24780 39090 24900 39210
rect 25500 39090 25620 39210
rect 26460 39090 26580 39210
rect 26940 39090 27060 39210
rect 27900 39090 28020 39210
rect 31020 39090 31140 39210
rect 32460 39090 32580 39210
rect 33420 39090 33540 39210
rect 34860 39090 34980 39210
rect 36060 39090 36180 39210
rect 36780 39090 36900 39210
rect 38220 39090 38340 39210
rect 38940 39090 39060 39210
rect 39660 39090 39780 39210
rect 40380 39090 40500 39210
rect 42060 39090 42180 39210
rect 43020 39090 43140 39210
rect 43740 39090 43860 39210
rect 44940 39090 45060 39210
rect 45900 39090 46020 39210
rect 46620 39090 46740 39210
rect 47580 39090 47700 39210
rect 48300 39090 48420 39210
rect 49740 39090 49860 39210
rect 6540 38790 6660 38910
rect 10620 38790 10740 38910
rect 15660 38790 15780 38910
rect 18780 38790 18900 38910
rect 23820 38790 23940 38910
rect 28140 38790 28260 38910
rect 41820 38790 41940 38910
rect 44700 38790 44820 38910
rect 7260 37290 7380 37410
rect 23820 37290 23940 37410
rect 31260 37290 31380 37410
rect 38940 37290 39060 37410
rect 41580 37290 41700 37410
rect 43740 37290 43860 37410
rect 6060 36990 6180 37110
rect 7020 36990 7140 37110
rect 8220 36990 8340 37110
rect 8940 36990 9060 37110
rect 10860 36990 10980 37110
rect 12060 36990 12180 37110
rect 12780 36990 12900 37110
rect 14940 36990 15060 37110
rect 15660 36990 15780 37110
rect 17340 36990 17460 37110
rect 18060 36990 18180 37110
rect 19500 36990 19620 37110
rect 20940 36990 21060 37110
rect 22380 36990 22500 37110
rect 24060 36990 24180 37110
rect 25500 36990 25620 37110
rect 26460 36990 26580 37110
rect 27180 36990 27300 37110
rect 27900 36990 28020 37110
rect 29100 36990 29220 37110
rect 30060 36990 30180 37110
rect 30780 36990 30900 37110
rect 31500 36990 31620 37110
rect 31980 36990 32100 37110
rect 32700 36990 32820 37110
rect 33660 36990 33780 37110
rect 34620 36990 34740 37110
rect 35580 36990 35700 37110
rect 37020 36990 37140 37110
rect 39180 36990 39300 37110
rect 40140 36990 40260 37110
rect 40620 36990 40740 37110
rect 41820 36990 41940 37110
rect 42300 36990 42420 37110
rect 43020 36990 43140 37110
rect 43500 36990 43620 37110
rect 44460 36990 44580 37110
rect 45180 36990 45300 37110
rect 46140 36990 46260 37110
rect 47580 36990 47700 37110
rect 48300 36990 48420 37110
rect 49740 36990 49860 37110
rect 5820 36690 5940 36810
rect 8700 36690 8820 36810
rect 11100 36690 11220 36810
rect 12540 36690 12660 36810
rect 15420 36690 15540 36810
rect 18300 36690 18420 36810
rect 19740 36690 19860 36810
rect 21180 36690 21300 36810
rect 22620 36690 22740 36810
rect 25260 36690 25380 36810
rect 26700 36690 26820 36810
rect 28140 36690 28260 36810
rect 29340 36690 29460 36810
rect 30300 36690 30420 36810
rect 32460 36690 32580 36810
rect 33420 36690 33540 36810
rect 34860 36690 34980 36810
rect 36300 36690 36420 36810
rect 39900 36690 40020 36810
rect 40380 36690 40500 36810
rect 40860 36690 40980 36810
rect 42780 36690 42900 36810
rect 44700 36690 44820 36810
rect 46380 36690 46500 36810
rect 47820 36690 47940 36810
rect 49500 36690 49620 36810
rect 5580 36390 5700 36510
rect 8220 36390 8340 36510
rect 11340 36390 11460 36510
rect 12060 36390 12180 36510
rect 14940 36390 15060 36510
rect 17100 36390 17220 36510
rect 18540 36390 18660 36510
rect 19980 36390 20100 36510
rect 21420 36390 21540 36510
rect 22860 36390 22980 36510
rect 25020 36390 25140 36510
rect 27180 36390 27300 36510
rect 28380 36390 28500 36510
rect 29580 36390 29700 36510
rect 30780 36390 30900 36510
rect 31980 36390 32100 36510
rect 33180 36390 33300 36510
rect 35100 36390 35220 36510
rect 42300 36390 42420 36510
rect 45180 36390 45300 36510
rect 46620 36390 46740 36510
rect 48300 36390 48420 36510
rect 49260 36390 49380 36510
rect 16620 36090 16740 36210
rect 20700 33990 20820 34110
rect 6540 33690 6660 33810
rect 7740 33690 7860 33810
rect 15660 33690 15780 33810
rect 17340 33690 17460 33810
rect 19260 33690 19380 33810
rect 21180 33690 21300 33810
rect 24060 33690 24180 33810
rect 25500 33690 25620 33810
rect 31020 33690 31140 33810
rect 32700 33690 32820 33810
rect 33660 33690 33780 33810
rect 35100 33690 35220 33810
rect 36540 33690 36660 33810
rect 37500 33690 37620 33810
rect 39420 33690 39540 33810
rect 40860 33690 40980 33810
rect 42060 33690 42180 33810
rect 43740 33690 43860 33810
rect 46860 33690 46980 33810
rect 47580 33690 47700 33810
rect 49020 33690 49140 33810
rect 7020 33390 7140 33510
rect 8220 33390 8340 33510
rect 9900 33390 10020 33510
rect 12060 33390 12180 33510
rect 15420 33390 15540 33510
rect 16860 33390 16980 33510
rect 19500 33390 19620 33510
rect 23580 33390 23700 33510
rect 25020 33390 25140 33510
rect 26700 33390 26820 33510
rect 31260 33390 31380 33510
rect 32220 33390 32340 33510
rect 33420 33390 33540 33510
rect 34860 33390 34980 33510
rect 36300 33390 36420 33510
rect 37740 33390 37860 33510
rect 39180 33390 39300 33510
rect 40380 33390 40500 33510
rect 41820 33390 41940 33510
rect 43260 33390 43380 33510
rect 44940 33390 45060 33510
rect 46380 33390 46500 33510
rect 47820 33390 47940 33510
rect 49260 33390 49380 33510
rect 6540 33090 6660 33210
rect 7260 33090 7380 33210
rect 7740 33090 7860 33210
rect 8460 33090 8580 33210
rect 8940 33090 9060 33210
rect 10380 33090 10500 33210
rect 11100 33090 11220 33210
rect 12540 33090 12660 33210
rect 13740 33090 13860 33210
rect 15180 33090 15300 33210
rect 16620 33090 16740 33210
rect 17340 33090 17460 33210
rect 19740 33090 19860 33210
rect 21420 33090 21540 33210
rect 23340 33090 23460 33210
rect 24060 33090 24180 33210
rect 24780 33090 24900 33210
rect 25500 33090 25620 33210
rect 25980 33090 26100 33210
rect 27420 33090 27540 33210
rect 30300 33090 30420 33210
rect 31500 33090 31620 33210
rect 31980 33090 32100 33210
rect 32700 33090 32820 33210
rect 33180 33090 33300 33210
rect 34620 33090 34740 33210
rect 36060 33090 36180 33210
rect 37980 33090 38100 33210
rect 38940 33090 39060 33210
rect 40140 33090 40260 33210
rect 40860 33090 40980 33210
rect 41580 33090 41700 33210
rect 43020 33090 43140 33210
rect 43740 33090 43860 33210
rect 44220 33090 44340 33210
rect 45660 33090 45780 33210
rect 46140 33090 46260 33210
rect 46860 33090 46980 33210
rect 48060 33090 48180 33210
rect 49500 33090 49620 33210
rect 13980 32790 14100 32910
rect 30540 32790 30660 32910
rect 24060 31290 24180 31410
rect 27420 31290 27540 31410
rect 28620 31290 28740 31410
rect 40860 31290 40980 31410
rect 5340 30990 5460 31110
rect 6780 30990 6900 31110
rect 7980 30990 8100 31110
rect 8700 30990 8820 31110
rect 10140 30990 10260 31110
rect 11100 30990 11220 31110
rect 12540 30990 12660 31110
rect 14700 30990 14820 31110
rect 16140 30990 16260 31110
rect 17100 30990 17220 31110
rect 18540 30990 18660 31110
rect 19260 30990 19380 31110
rect 20700 30990 20820 31110
rect 21180 30990 21300 31110
rect 22140 30990 22260 31110
rect 22860 30990 22980 31110
rect 23820 30990 23940 31110
rect 25500 30990 25620 31110
rect 25980 30990 26100 31110
rect 26700 30990 26820 31110
rect 27180 30990 27300 31110
rect 28140 30990 28260 31110
rect 28860 30990 28980 31110
rect 29100 30990 29220 31110
rect 29820 30990 29940 31110
rect 30780 30990 30900 31110
rect 32220 30990 32340 31110
rect 33180 30990 33300 31110
rect 34620 30990 34740 31110
rect 36060 30990 36180 31110
rect 36780 30990 36900 31110
rect 37740 30990 37860 31110
rect 38940 30990 39060 31110
rect 39660 30990 39780 31110
rect 40620 30990 40740 31110
rect 42060 30990 42180 31110
rect 43020 30990 43140 31110
rect 43740 30990 43860 31110
rect 44460 30990 44580 31110
rect 45180 30990 45300 31110
rect 46620 30990 46740 31110
rect 48060 30990 48180 31110
rect 49500 30990 49620 31110
rect 5820 30690 5940 30810
rect 8220 30690 8340 30810
rect 9900 30690 10020 30810
rect 11820 30690 11940 30810
rect 15660 30690 15780 30810
rect 18060 30690 18180 30810
rect 19980 30690 20100 30810
rect 21420 30690 21540 30810
rect 22620 30690 22740 30810
rect 26460 30690 26580 30810
rect 27900 30690 28020 30810
rect 29580 30690 29700 30810
rect 31500 30690 31620 30810
rect 33420 30690 33540 30810
rect 34860 30690 34980 30810
rect 36540 30690 36660 30810
rect 37980 30690 38100 30810
rect 39180 30690 39300 30810
rect 41820 30690 41940 30810
rect 43500 30690 43620 30810
rect 44700 30690 44820 30810
rect 46380 30690 46500 30810
rect 48780 30690 48900 30810
rect 8700 30390 8820 30510
rect 9660 30390 9780 30510
rect 21660 30390 21780 30510
rect 22140 30390 22260 30510
rect 25260 30390 25380 30510
rect 25980 30390 26100 30510
rect 27660 30390 27780 30510
rect 29100 30390 29220 30510
rect 33660 30390 33780 30510
rect 35100 30390 35220 30510
rect 36060 30390 36180 30510
rect 38220 30390 38340 30510
rect 39660 30390 39780 30510
rect 41580 30390 41700 30510
rect 43020 30390 43140 30510
rect 45180 30390 45300 30510
rect 46140 30390 46260 30510
rect 24780 30090 24900 30210
rect 13740 27990 13860 28110
rect 9180 27690 9300 27810
rect 11820 27690 11940 27810
rect 12540 27690 12660 27810
rect 13260 27690 13380 27810
rect 14220 27690 14340 27810
rect 15900 27690 16020 27810
rect 16620 27690 16740 27810
rect 18540 27690 18660 27810
rect 19260 27690 19380 27810
rect 21420 27690 21540 27810
rect 22620 27690 22740 27810
rect 24060 27690 24180 27810
rect 25500 27690 25620 27810
rect 26940 27690 27060 27810
rect 28380 27690 28500 27810
rect 30300 27690 30420 27810
rect 31740 27690 31860 27810
rect 35340 27690 35460 27810
rect 36540 27690 36660 27810
rect 37500 27690 37620 27810
rect 39180 27690 39300 27810
rect 42060 27690 42180 27810
rect 43020 27690 43140 27810
rect 45180 27690 45300 27810
rect 46620 27690 46740 27810
rect 49020 27690 49140 27810
rect 49980 27690 50100 27810
rect 7740 27390 7860 27510
rect 8940 27390 9060 27510
rect 9900 27390 10020 27510
rect 11340 27390 11460 27510
rect 12300 27390 12420 27510
rect 13020 27390 13140 27510
rect 15660 27390 15780 27510
rect 16860 27390 16980 27510
rect 18300 27390 18420 27510
rect 19740 27390 19860 27510
rect 21180 27390 21300 27510
rect 22380 27390 22500 27510
rect 23820 27390 23940 27510
rect 25260 27390 25380 27510
rect 26700 27390 26820 27510
rect 28860 27390 28980 27510
rect 30540 27390 30660 27510
rect 32220 27390 32340 27510
rect 33660 27390 33780 27510
rect 35100 27390 35220 27510
rect 36300 27390 36420 27510
rect 37740 27390 37860 27510
rect 38940 27390 39060 27510
rect 40380 27390 40500 27510
rect 41820 27390 41940 27510
rect 43500 27390 43620 27510
rect 44700 27390 44820 27510
rect 46140 27390 46260 27510
rect 47340 27390 47460 27510
rect 47820 27390 47940 27510
rect 48300 27390 48420 27510
rect 48780 27390 48900 27510
rect 49500 27390 49620 27510
rect 7020 27090 7140 27210
rect 8460 27090 8580 27210
rect 8700 27090 8820 27210
rect 9420 27090 9540 27210
rect 10860 27090 10980 27210
rect 11100 27090 11220 27210
rect 11820 27090 11940 27210
rect 12060 27090 12180 27210
rect 12780 27090 12900 27210
rect 14460 27090 14580 27210
rect 15420 27090 15540 27210
rect 17100 27090 17220 27210
rect 18060 27090 18180 27210
rect 19260 27090 19380 27210
rect 19980 27090 20100 27210
rect 20940 27090 21060 27210
rect 22140 27090 22260 27210
rect 23580 27090 23700 27210
rect 25020 27090 25140 27210
rect 26460 27090 26580 27210
rect 28380 27090 28500 27210
rect 29100 27090 29220 27210
rect 30780 27090 30900 27210
rect 31740 27090 31860 27210
rect 32460 27090 32580 27210
rect 32940 27090 33060 27210
rect 34380 27090 34500 27210
rect 34860 27090 34980 27210
rect 36060 27090 36180 27210
rect 37980 27090 38100 27210
rect 38700 27090 38820 27210
rect 39660 27090 39780 27210
rect 41100 27090 41220 27210
rect 41580 27090 41700 27210
rect 43020 27090 43140 27210
rect 43740 27090 43860 27210
rect 44460 27090 44580 27210
rect 45180 27090 45300 27210
rect 45900 27090 46020 27210
rect 46620 27090 46740 27210
rect 47100 27090 47220 27210
rect 47580 27090 47700 27210
rect 48060 27090 48180 27210
rect 48540 27090 48660 27210
rect 49260 27090 49380 27210
rect 49980 27090 50100 27210
rect 46860 26790 46980 26910
rect 12060 25290 12180 25410
rect 13980 25290 14100 25410
rect 30540 25290 30660 25410
rect 32460 25290 32580 25410
rect 43260 25290 43380 25410
rect 44460 25290 44580 25410
rect 5340 24990 5460 25110
rect 6780 24990 6900 25110
rect 7020 24990 7140 25110
rect 7740 24990 7860 25110
rect 8460 24990 8580 25110
rect 8700 24990 8820 25110
rect 9420 24990 9540 25110
rect 10860 24990 10980 25110
rect 12540 24990 12660 25110
rect 13740 24990 13860 25110
rect 14940 24990 15060 25110
rect 15660 24990 15780 25110
rect 21180 24990 21300 25110
rect 23100 24990 23220 25110
rect 25500 24990 25620 25110
rect 26940 24990 27060 25110
rect 27900 24990 28020 25110
rect 28620 24990 28740 25110
rect 30300 24990 30420 25110
rect 31020 24990 31140 25110
rect 31740 24990 31860 25110
rect 32220 24990 32340 25110
rect 33180 24990 33300 25110
rect 34620 24990 34740 25110
rect 36060 24990 36180 25110
rect 37500 24990 37620 25110
rect 38940 24990 39060 25110
rect 40380 24990 40500 25110
rect 41820 24990 41940 25110
rect 43500 24990 43620 25110
rect 44700 24990 44820 25110
rect 47820 24990 47940 25110
rect 49260 24990 49380 25110
rect 6060 24690 6180 24810
rect 7260 24690 7380 24810
rect 8220 24690 8340 24810
rect 8940 24690 9060 24810
rect 10140 24690 10260 24810
rect 12060 24690 12180 24810
rect 12780 24690 12900 24810
rect 15420 24690 15540 24810
rect 20940 24690 21060 24810
rect 23340 24690 23460 24810
rect 26220 24690 26340 24810
rect 28380 24690 28500 24810
rect 31500 24690 31620 24810
rect 33420 24690 33540 24810
rect 34860 24690 34980 24810
rect 36300 24690 36420 24810
rect 37740 24690 37860 24810
rect 39180 24690 39300 24810
rect 40620 24690 40740 24810
rect 42060 24690 42180 24810
rect 43740 24690 43860 24810
rect 48540 24690 48660 24810
rect 7500 24390 7620 24510
rect 7740 24390 7860 24510
rect 9180 24390 9300 24510
rect 14940 24390 15060 24510
rect 20700 24390 20820 24510
rect 23580 24390 23700 24510
rect 27900 24390 28020 24510
rect 31020 24390 31140 24510
rect 33660 24390 33780 24510
rect 35100 24390 35220 24510
rect 36540 24390 36660 24510
rect 37980 24390 38100 24510
rect 39420 24390 39540 24510
rect 40860 24390 40980 24510
rect 42300 24390 42420 24510
rect 8700 21690 8820 21810
rect 10140 21690 10260 21810
rect 11100 21690 11220 21810
rect 18540 21690 18660 21810
rect 22140 21690 22260 21810
rect 26220 21690 26340 21810
rect 27900 21690 28020 21810
rect 29580 21690 29700 21810
rect 31020 21690 31140 21810
rect 32460 21690 32580 21810
rect 33660 21690 33780 21810
rect 35100 21690 35220 21810
rect 36300 21690 36420 21810
rect 38940 21690 39060 21810
rect 40860 21690 40980 21810
rect 41580 21690 41700 21810
rect 6060 21390 6180 21510
rect 8460 21390 8580 21510
rect 9900 21390 10020 21510
rect 11580 21390 11700 21510
rect 14940 21390 15060 21510
rect 18300 21390 18420 21510
rect 19500 21390 19620 21510
rect 21180 21390 21300 21510
rect 22620 21390 22740 21510
rect 26700 21390 26820 21510
rect 28380 21390 28500 21510
rect 29340 21390 29460 21510
rect 30540 21390 30660 21510
rect 32220 21390 32340 21510
rect 33420 21390 33540 21510
rect 34860 21390 34980 21510
rect 36060 21390 36180 21510
rect 37500 21390 37620 21510
rect 39420 21390 39540 21510
rect 40620 21390 40740 21510
rect 42060 21390 42180 21510
rect 43740 21390 43860 21510
rect 44940 21390 45060 21510
rect 46620 21390 46740 21510
rect 48780 21390 48900 21510
rect 49260 21390 49380 21510
rect 49740 21390 49860 21510
rect 5340 21090 5460 21210
rect 6780 21090 6900 21210
rect 8220 21090 8340 21210
rect 9660 21090 9780 21210
rect 11100 21090 11220 21210
rect 11820 21090 11940 21210
rect 14220 21090 14340 21210
rect 15660 21090 15780 21210
rect 16860 21090 16980 21210
rect 18060 21090 18180 21210
rect 18780 21090 18900 21210
rect 20220 21090 20340 21210
rect 20460 21090 20580 21210
rect 21900 21090 22020 21210
rect 22140 21090 22260 21210
rect 22860 21090 22980 21210
rect 25260 21090 25380 21210
rect 26220 21090 26340 21210
rect 26940 21090 27060 21210
rect 27900 21090 28020 21210
rect 28620 21090 28740 21210
rect 29100 21090 29220 21210
rect 30300 21090 30420 21210
rect 31020 21090 31140 21210
rect 31980 21090 32100 21210
rect 33180 21090 33300 21210
rect 34620 21090 34740 21210
rect 35820 21090 35940 21210
rect 36780 21090 36900 21210
rect 38220 21090 38340 21210
rect 38940 21090 39060 21210
rect 39660 21090 39780 21210
rect 40380 21090 40500 21210
rect 41580 21090 41700 21210
rect 42300 21090 42420 21210
rect 43500 21090 43620 21210
rect 44220 21090 44340 21210
rect 45660 21090 45780 21210
rect 45900 21090 46020 21210
rect 47340 21090 47460 21210
rect 47820 21090 47940 21210
rect 49020 21090 49140 21210
rect 49500 21090 49620 21210
rect 17100 20790 17220 20910
rect 25020 20790 25140 20910
rect 43260 20790 43380 20910
rect 47580 20790 47700 20910
rect 16140 19290 16260 19410
rect 27420 19290 27540 19410
rect 36780 19290 36900 19410
rect 41580 19290 41700 19410
rect 47580 19290 47700 19410
rect 5580 18990 5700 19110
rect 6300 18990 6420 19110
rect 8940 18990 9060 19110
rect 10380 18990 10500 19110
rect 11580 18990 11700 19110
rect 13020 18990 13140 19110
rect 13500 18990 13620 19110
rect 14940 18990 15060 19110
rect 15660 18990 15780 19110
rect 17820 18990 17940 19110
rect 18540 18990 18660 19110
rect 19500 18990 19620 19110
rect 20940 18990 21060 19110
rect 22140 18990 22260 19110
rect 23580 18990 23700 19110
rect 24540 18990 24660 19110
rect 25980 18990 26100 19110
rect 26220 18990 26340 19110
rect 26940 18990 27060 19110
rect 27180 18990 27300 19110
rect 28380 18990 28500 19110
rect 29100 18990 29220 19110
rect 30540 18990 30660 19110
rect 31980 18990 32100 19110
rect 33180 18990 33300 19110
rect 33900 18990 34020 19110
rect 35820 18990 35940 19110
rect 37260 18990 37380 19110
rect 37980 18990 38100 19110
rect 38940 18990 39060 19110
rect 40380 18990 40500 19110
rect 41820 18990 41940 19110
rect 43020 18990 43140 19110
rect 43500 18990 43620 19110
rect 44460 18990 44580 19110
rect 45180 18990 45300 19110
rect 46140 18990 46260 19110
rect 47820 18990 47940 19110
rect 49020 18990 49140 19110
rect 49740 18990 49860 19110
rect 6060 18690 6180 18810
rect 9660 18690 9780 18810
rect 12540 18690 12660 18810
rect 14220 18690 14340 18810
rect 15420 18690 15540 18810
rect 16140 18690 16260 18810
rect 18300 18690 18420 18810
rect 19740 18690 19860 18810
rect 21180 18690 21300 18810
rect 22380 18690 22500 18810
rect 23820 18690 23940 18810
rect 25260 18690 25380 18810
rect 26460 18690 26580 18810
rect 28860 18690 28980 18810
rect 30780 18690 30900 18810
rect 32220 18690 32340 18810
rect 33420 18690 33540 18810
rect 36060 18690 36180 18810
rect 36780 18690 36900 18810
rect 37500 18690 37620 18810
rect 38220 18690 38340 18810
rect 39180 18690 39300 18810
rect 40620 18690 40740 18810
rect 42780 18690 42900 18810
rect 43260 18690 43380 18810
rect 43740 18690 43860 18810
rect 44700 18690 44820 18810
rect 46380 18690 46500 18810
rect 48060 18690 48180 18810
rect 49260 18690 49380 18810
rect 5580 18390 5700 18510
rect 17820 18390 17940 18510
rect 19980 18390 20100 18510
rect 21420 18390 21540 18510
rect 22620 18390 22740 18510
rect 24060 18390 24180 18510
rect 26940 18390 27060 18510
rect 28380 18390 28500 18510
rect 31020 18390 31140 18510
rect 32460 18390 32580 18510
rect 33900 18390 34020 18510
rect 36300 18390 36420 18510
rect 38460 18390 38580 18510
rect 39420 18390 39540 18510
rect 40860 18390 40980 18510
rect 45180 18390 45300 18510
rect 46620 18390 46740 18510
rect 49740 18390 49860 18510
rect 6780 15690 6900 15810
rect 18060 15690 18180 15810
rect 19740 15690 19860 15810
rect 21420 15690 21540 15810
rect 22140 15690 22260 15810
rect 24060 15690 24180 15810
rect 24780 15690 24900 15810
rect 28380 15690 28500 15810
rect 29580 15690 29700 15810
rect 32220 15690 32340 15810
rect 33660 15690 33780 15810
rect 35100 15690 35220 15810
rect 36780 15690 36900 15810
rect 38220 15690 38340 15810
rect 45180 15690 45300 15810
rect 46620 15690 46740 15810
rect 47580 15690 47700 15810
rect 49740 15690 49860 15810
rect 6540 15390 6660 15510
rect 8460 15390 8580 15510
rect 10140 15390 10260 15510
rect 12060 15390 12180 15510
rect 14220 15390 14340 15510
rect 15660 15390 15780 15510
rect 16620 15390 16740 15510
rect 17340 15390 17460 15510
rect 18540 15390 18660 15510
rect 19500 15390 19620 15510
rect 20940 15390 21060 15510
rect 22620 15390 22740 15510
rect 23820 15390 23940 15510
rect 25020 15390 25140 15510
rect 26460 15390 26580 15510
rect 28140 15390 28260 15510
rect 29340 15390 29460 15510
rect 31020 15390 31140 15510
rect 32460 15390 32580 15510
rect 33420 15390 33540 15510
rect 34860 15390 34980 15510
rect 36300 15390 36420 15510
rect 37980 15390 38100 15510
rect 39420 15390 39540 15510
rect 42300 15390 42420 15510
rect 44700 15390 44820 15510
rect 46380 15390 46500 15510
rect 47820 15390 47940 15510
rect 49260 15390 49380 15510
rect 6300 15090 6420 15210
rect 7740 15090 7860 15210
rect 9180 15090 9300 15210
rect 9420 15090 9540 15210
rect 10860 15090 10980 15210
rect 11100 15090 11220 15210
rect 12540 15090 12660 15210
rect 13260 15090 13380 15210
rect 14700 15090 14820 15210
rect 14940 15090 15060 15210
rect 16380 15090 16500 15210
rect 16860 15090 16980 15210
rect 17580 15090 17700 15210
rect 18060 15090 18180 15210
rect 18780 15090 18900 15210
rect 19260 15090 19380 15210
rect 20700 15090 20820 15210
rect 21420 15090 21540 15210
rect 22140 15090 22260 15210
rect 22860 15090 22980 15210
rect 23580 15090 23700 15210
rect 25260 15090 25380 15210
rect 25740 15090 25860 15210
rect 27180 15090 27300 15210
rect 27900 15090 28020 15210
rect 29100 15090 29220 15210
rect 30300 15090 30420 15210
rect 31740 15090 31860 15210
rect 32700 15090 32820 15210
rect 33180 15090 33300 15210
rect 34620 15090 34740 15210
rect 36060 15090 36180 15210
rect 36780 15090 36900 15210
rect 37740 15090 37860 15210
rect 38700 15090 38820 15210
rect 40140 15090 40260 15210
rect 41580 15090 41700 15210
rect 43020 15090 43140 15210
rect 44460 15090 44580 15210
rect 45180 15090 45300 15210
rect 46140 15090 46260 15210
rect 48060 15090 48180 15210
rect 49020 15090 49140 15210
rect 49740 15090 49860 15210
rect 17340 14790 17460 14910
rect 17820 14790 17940 14910
rect 7260 12990 7380 13110
rect 8940 12990 9060 13110
rect 9420 12990 9540 13110
rect 9900 12990 10020 13110
rect 10860 12990 10980 13110
rect 12060 12990 12180 13110
rect 12780 12990 12900 13110
rect 15900 12990 16020 13110
rect 16620 12990 16740 13110
rect 17340 12990 17460 13110
rect 17580 12990 17700 13110
rect 19020 12990 19140 13110
rect 19260 12990 19380 13110
rect 20700 12990 20820 13110
rect 21900 12990 22020 13110
rect 23340 12990 23460 13110
rect 25020 12990 25140 13110
rect 25740 12990 25860 13110
rect 26700 12990 26820 13110
rect 29100 12990 29220 13110
rect 29820 12990 29940 13110
rect 30300 12990 30420 13110
rect 31020 12990 31140 13110
rect 32460 12990 32580 13110
rect 32940 12990 33060 13110
rect 34380 12990 34500 13110
rect 34620 12990 34740 13110
rect 35340 12990 35460 13110
rect 36060 12990 36180 13110
rect 37500 12990 37620 13110
rect 38940 12990 39060 13110
rect 40140 12990 40260 13110
rect 40860 12990 40980 13110
rect 41580 12990 41700 13110
rect 43260 12990 43380 13110
rect 44460 12990 44580 13110
rect 45180 12990 45300 13110
rect 46140 12990 46260 13110
rect 47580 12990 47700 13110
rect 48300 12990 48420 13110
rect 49740 12990 49860 13110
rect 7020 12690 7140 12810
rect 9180 12690 9300 12810
rect 9660 12690 9780 12810
rect 11100 12690 11220 12810
rect 12540 12690 12660 12810
rect 16140 12690 16260 12810
rect 17100 12690 17220 12810
rect 18300 12690 18420 12810
rect 19740 12690 19860 12810
rect 22860 12690 22980 12810
rect 25260 12690 25380 12810
rect 26940 12690 27060 12810
rect 29340 12690 29460 12810
rect 30780 12690 30900 12810
rect 32220 12690 32340 12810
rect 33660 12690 33780 12810
rect 34860 12690 34980 12810
rect 36300 12690 36420 12810
rect 37740 12690 37860 12810
rect 39180 12690 39300 12810
rect 40620 12690 40740 12810
rect 43500 12690 43620 12810
rect 44700 12690 44820 12810
rect 46380 12690 46500 12810
rect 47820 12690 47940 12810
rect 49500 12690 49620 12810
rect 6780 12390 6900 12510
rect 11340 12390 11460 12510
rect 12060 12390 12180 12510
rect 16380 12390 16500 12510
rect 16620 12390 16740 12510
rect 25740 12390 25860 12510
rect 27180 12390 27300 12510
rect 29820 12390 29940 12510
rect 30300 12390 30420 12510
rect 31980 12390 32100 12510
rect 35340 12390 35460 12510
rect 36540 12390 36660 12510
rect 37980 12390 38100 12510
rect 39420 12390 39540 12510
rect 40140 12390 40260 12510
rect 41820 12390 41940 12510
rect 43740 12390 43860 12510
rect 45180 12390 45300 12510
rect 46620 12390 46740 12510
rect 48300 12390 48420 12510
rect 49260 12390 49380 12510
rect 42300 12090 42420 12210
rect 9660 9990 9780 10110
rect 35580 9990 35700 10110
rect 37740 9990 37860 10110
rect 5580 9690 5700 9810
rect 7260 9690 7380 9810
rect 10140 9690 10260 9810
rect 11340 9690 11460 9810
rect 16860 9690 16980 9810
rect 21180 9690 21300 9810
rect 24300 9690 24420 9810
rect 28380 9690 28500 9810
rect 32460 9690 32580 9810
rect 36060 9690 36180 9810
rect 37260 9690 37380 9810
rect 38220 9690 38340 9810
rect 39660 9690 39780 9810
rect 40860 9690 40980 9810
rect 42060 9690 42180 9810
rect 47580 9690 47700 9810
rect 49020 9690 49140 9810
rect 6060 9390 6180 9510
rect 7020 9390 7140 9510
rect 8460 9390 8580 9510
rect 11580 9390 11700 9510
rect 14460 9390 14580 9510
rect 16620 9390 16740 9510
rect 18300 9390 18420 9510
rect 19980 9390 20100 9510
rect 21420 9390 21540 9510
rect 22620 9390 22740 9510
rect 24060 9390 24180 9510
rect 26220 9390 26340 9510
rect 28140 9390 28260 9510
rect 31980 9390 32100 9510
rect 33660 9390 33780 9510
rect 37020 9390 37140 9510
rect 39180 9390 39300 9510
rect 40620 9390 40740 9510
rect 41820 9390 41940 9510
rect 43260 9390 43380 9510
rect 45900 9390 46020 9510
rect 47820 9390 47940 9510
rect 49260 9390 49380 9510
rect 5580 9090 5700 9210
rect 6300 9090 6420 9210
rect 6780 9090 6900 9210
rect 7740 9090 7860 9210
rect 9180 9090 9300 9210
rect 10380 9090 10500 9210
rect 11820 9090 11940 9210
rect 13740 9090 13860 9210
rect 15180 9090 15300 9210
rect 16380 9090 16500 9210
rect 17340 9090 17460 9210
rect 18780 9090 18900 9210
rect 19260 9090 19380 9210
rect 20700 9090 20820 9210
rect 21660 9090 21780 9210
rect 21900 9090 22020 9210
rect 23340 9090 23460 9210
rect 23820 9090 23940 9210
rect 25500 9090 25620 9210
rect 26940 9090 27060 9210
rect 27900 9090 28020 9210
rect 29340 9090 29460 9210
rect 30780 9090 30900 9210
rect 31740 9090 31860 9210
rect 32460 9090 32580 9210
rect 33180 9090 33300 9210
rect 34620 9090 34740 9210
rect 36300 9090 36420 9210
rect 36780 9090 36900 9210
rect 38460 9090 38580 9210
rect 38940 9090 39060 9210
rect 39660 9090 39780 9210
rect 40380 9090 40500 9210
rect 41580 9090 41700 9210
rect 42540 9090 42660 9210
rect 43980 9090 44100 9210
rect 45180 9090 45300 9210
rect 46620 9090 46740 9210
rect 48060 9090 48180 9210
rect 49500 9090 49620 9210
rect 29580 8790 29700 8910
rect 30540 8790 30660 8910
rect 8220 7290 8340 7410
rect 14460 7290 14580 7410
rect 15420 7290 15540 7410
rect 18060 7290 18180 7410
rect 43260 7290 43380 7410
rect 46620 7290 46740 7410
rect 5580 6990 5700 7110
rect 7020 6990 7140 7110
rect 7980 6990 8100 7110
rect 8700 6990 8820 7110
rect 9420 6990 9540 7110
rect 9900 6990 10020 7110
rect 10860 6990 10980 7110
rect 11580 6990 11700 7110
rect 12300 6990 12420 7110
rect 13980 6990 14100 7110
rect 15660 6990 15780 7110
rect 18300 6990 18420 7110
rect 20700 6990 20820 7110
rect 23340 6990 23460 7110
rect 25740 6990 25860 7110
rect 27180 6990 27300 7110
rect 27900 6990 28020 7110
rect 29100 6990 29220 7110
rect 30060 6990 30180 7110
rect 31500 6990 31620 7110
rect 31980 6990 32100 7110
rect 32700 6990 32820 7110
rect 33180 6990 33300 7110
rect 35100 6990 35220 7110
rect 36060 6990 36180 7110
rect 37500 6990 37620 7110
rect 38220 6990 38340 7110
rect 38940 6990 39060 7110
rect 40380 6990 40500 7110
rect 43500 6990 43620 7110
rect 44700 6990 44820 7110
rect 45180 6990 45300 7110
rect 46380 6990 46500 7110
rect 47340 6990 47460 7110
rect 48060 6990 48180 7110
rect 6300 6690 6420 6810
rect 9180 6690 9300 6810
rect 10140 6690 10260 6810
rect 11340 6690 11460 6810
rect 12540 6690 12660 6810
rect 13740 6690 13860 6810
rect 14460 6690 14580 6810
rect 15900 6690 16020 6810
rect 18540 6690 18660 6810
rect 20940 6690 21060 6810
rect 23580 6690 23700 6810
rect 26700 6690 26820 6810
rect 28140 6690 28260 6810
rect 29340 6690 29460 6810
rect 30780 6690 30900 6810
rect 32220 6690 32340 6810
rect 33420 6690 33540 6810
rect 34860 6690 34980 6810
rect 36300 6690 36420 6810
rect 37980 6690 38100 6810
rect 39180 6690 39300 6810
rect 40620 6690 40740 6810
rect 43740 6690 43860 6810
rect 44460 6690 44580 6810
rect 44940 6690 45060 6810
rect 45420 6690 45540 6810
rect 47820 6690 47940 6810
rect 8700 6390 8820 6510
rect 10380 6390 10500 6510
rect 10860 6390 10980 6510
rect 12780 6390 12900 6510
rect 21180 6390 21300 6510
rect 23820 6390 23940 6510
rect 28380 6390 28500 6510
rect 29580 6390 29700 6510
rect 32700 6390 32820 6510
rect 33660 6390 33780 6510
rect 34620 6390 34740 6510
rect 36540 6390 36660 6510
rect 37500 6390 37620 6510
rect 39420 6390 39540 6510
rect 40860 6390 40980 6510
rect 47340 6390 47460 6510
<< labels >>
rlabel metal3 60 43500 60 43500 6 P_15_
rlabel metal3 60 38100 60 38100 6 P_14_
rlabel metal3 60 32700 60 32700 6 P_13_
rlabel metal3 60 27300 60 27300 6 P_12_
rlabel metal3 60 21900 60 21900 6 P_11_
rlabel metal3 60 16500 60 16500 6 P_10_
rlabel metal3 60 11100 60 11100 6 P_9_
rlabel metal3 60 5700 60 5700 6 P_8_
rlabel metal2 45720 49140 45720 49140 6 P_5_
rlabel metal2 36600 49140 36600 49140 6 P_4_
rlabel metal2 27720 49140 27720 49140 6 P_3_
rlabel metal2 18600 49140 18600 49140 6 P_2_
rlabel metal2 9480 49140 9480 49140 6 P_1_
rlabel metal2 36600 30 36600 30 6 A_7_
rlabel metal2 30600 30 30600 30 6 A_6_
rlabel metal2 24600 30 24600 30 6 A_5_
rlabel metal2 18600 30 18600 30 6 A_4_
rlabel metal2 12600 30 12600 30 6 A_3_
rlabel metal2 6600 30 6600 30 6 A_2_
rlabel metal3 55260 36600 55260 36600 6 B_6_
rlabel metal3 55260 24600 55260 24600 6 B_5_
rlabel metal3 55260 12600 55260 12600 6 B_4_
rlabel metal2 48600 30 48600 30 6 B_1_
rlabel metal2 42600 30 42600 30 6 B_0_
rlabel metal2 14520 49140 14520 49140 6 P_0_
rlabel metal3 55260 46950 55260 46950 6 B_7_
rlabel metal3 60 780 60 780 6 P_7_
rlabel metal3 55260 1080 55260 1080 6 B_3_
rlabel metal2 40410 30 40410 30 6 B_2_
rlabel metal2 53730 19830 53730 19830 6 vdd
rlabel metal1 37860 3450 37860 3450 6 gnd
rlabel metal3 60 46650 60 46650 6 A_0_
rlabel metal2 840 30 840 30 4 A_1_
rlabel metal2 54510 49140 54510 49140 4 P_6_
<< end >>

magic
tech scmos
timestamp 1053022145
<< nwell >>
rect -8 48 46 105
<< ntransistor >>
rect 9 6 11 26
rect 14 6 16 26
rect 26 6 28 26
rect 31 6 33 26
<< ptransistor >>
rect 7 54 9 94
rect 15 54 17 94
rect 23 54 25 94
rect 31 54 33 94
<< ndiffusion >>
rect 8 6 9 26
rect 11 6 14 26
rect 16 6 17 26
rect 25 6 26 26
rect 28 6 31 26
rect 33 6 34 26
<< pdiffusion >>
rect 6 57 7 94
rect 2 54 7 57
rect 9 60 10 94
rect 14 60 15 94
rect 9 54 15 60
rect 17 54 18 94
rect 22 54 23 94
rect 25 88 31 94
rect 25 54 26 88
rect 30 54 31 88
rect 33 54 34 94
<< ndcontact >>
rect 4 6 8 26
rect 17 6 25 26
rect 34 6 38 26
<< pdcontact >>
rect 2 57 6 94
rect 10 60 14 94
rect 18 54 22 94
rect 26 54 30 88
rect 34 54 38 94
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 31 94 33 96
rect 7 49 9 54
rect 15 53 17 54
rect 14 51 17 53
rect 4 29 6 47
rect 4 27 11 29
rect 9 26 11 27
rect 14 26 16 51
rect 23 40 25 54
rect 31 53 33 54
rect 31 51 35 53
rect 33 47 34 51
rect 24 39 25 40
rect 24 29 26 39
rect 33 31 35 47
rect 31 29 35 31
rect 24 27 28 29
rect 26 26 28 27
rect 31 26 33 29
rect 9 4 11 6
rect 14 4 16 6
rect 26 4 28 6
rect 31 4 33 6
<< polycontact >>
rect 6 45 10 49
rect 10 37 14 41
rect 34 47 38 51
rect 25 39 29 43
<< metal1 >>
rect -2 102 42 103
rect 2 98 14 102
rect 18 98 30 102
rect 34 98 42 102
rect -2 97 42 98
rect 10 94 14 97
rect 2 54 18 57
rect 22 91 34 94
rect 26 51 29 54
rect 2 45 6 47
rect 19 48 29 51
rect 19 47 22 48
rect 2 44 10 45
rect 2 43 6 44
rect 18 43 22 47
rect 34 43 38 47
rect 10 33 14 37
rect 19 26 22 43
rect 26 37 29 39
rect 26 33 30 37
rect 4 3 8 6
rect 34 3 38 6
rect -2 2 42 3
rect 2 -2 14 2
rect 18 -2 30 2
rect 34 -2 42 2
rect -2 -3 42 -2
<< m1p >>
rect 2 43 6 47
rect 18 43 22 47
rect 34 43 38 47
rect 10 33 14 37
rect 26 33 30 37
<< labels >>
rlabel metal1 4 0 4 0 1 gnd
rlabel metal1 4 100 4 100 5 vdd
rlabel metal1 36 45 36 45 1 C
rlabel metal1 28 35 28 35 1 D
rlabel metal1 20 45 20 45 1 Y
rlabel metal1 4 45 4 45 1 A
rlabel metal1 12 35 12 35 1 B
<< end >>

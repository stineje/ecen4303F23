magic
tech sky130A
magscale 1 2
timestamp 1606864426
<< checkpaint >>
rect -1269 2461 1546 2601
rect -1760 -1129 6260 2461
rect -1269 -1260 1546 -1129
<< nwell >>
rect -9 485 286 897
<< nmos >>
rect 80 115 110 219
rect 152 115 182 219
<< pmos >>
rect 80 521 110 773
rect 166 521 196 773
<< ndiff >>
rect 27 171 80 219
rect 27 131 35 171
rect 69 131 80 171
rect 27 115 80 131
rect 110 115 152 219
rect 182 171 235 219
rect 182 131 193 171
rect 227 131 235 171
rect 182 115 235 131
<< pdiff >>
rect 27 757 80 773
rect 27 697 35 757
rect 69 697 80 757
rect 27 521 80 697
rect 110 757 166 773
rect 110 561 121 757
rect 155 561 166 757
rect 110 521 166 561
rect 196 757 249 773
rect 196 629 207 757
rect 241 629 249 757
rect 196 521 249 629
<< ndiffc >>
rect 35 131 69 171
rect 193 131 227 171
<< pdiffc >>
rect 35 697 69 757
rect 121 561 155 757
rect 207 629 241 757
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 827 51 861
rect 85 827 109 861
rect 163 827 187 861
rect 221 827 245 861
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 827 85 861
rect 187 827 221 861
<< poly >>
rect 80 773 110 799
rect 166 773 196 799
rect 80 474 110 521
rect 37 458 110 474
rect 37 424 47 458
rect 81 424 110 458
rect 37 408 110 424
rect 80 219 110 408
rect 166 381 196 521
rect 152 365 210 381
rect 152 331 166 365
rect 200 331 210 365
rect 152 315 210 331
rect 152 219 182 315
rect 80 89 110 115
rect 152 89 182 115
<< polycont >>
rect 47 424 81 458
rect 166 331 200 365
<< locali >>
rect 0 867 286 888
rect 0 827 51 867
rect 85 827 187 867
rect 221 827 286 867
rect 35 757 69 827
rect 35 681 69 697
rect 121 757 155 773
rect 47 458 81 553
rect 47 408 81 424
rect 207 757 241 827
rect 207 613 241 629
rect 121 439 155 561
rect 195 365 229 479
rect 150 331 166 365
rect 200 331 229 365
rect 35 171 69 183
rect 35 115 69 131
rect 193 171 227 187
rect 193 61 227 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 286 61
rect 0 0 286 21
<< viali >>
rect 51 861 85 867
rect 51 833 85 861
rect 187 861 221 867
rect 187 833 221 861
rect 47 553 81 587
rect 121 405 155 439
rect 195 479 229 513
rect 35 183 69 217
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 867 286 888
rect 0 833 51 867
rect 85 833 187 867
rect 221 833 286 867
rect 0 827 286 833
rect 35 587 93 593
rect 35 553 47 587
rect 81 553 115 587
rect 35 547 93 553
rect 183 513 241 519
rect 161 479 195 513
rect 229 479 241 513
rect 183 473 241 479
rect 109 439 167 445
rect 109 405 121 439
rect 155 405 167 439
rect 109 399 167 405
rect 23 217 81 223
rect 121 217 155 399
rect 23 183 35 217
rect 69 183 155 217
rect 23 177 81 183
rect 0 55 286 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 286 55
rect 0 0 286 21
<< labels >>
rlabel metal1 136 374 136 374 1 Y
port 1 n
rlabel viali 64 570 64 570 1 A
port 2 n
rlabel viali 212 496 212 496 1 B
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 840 68 840 1 vdd
<< end >>

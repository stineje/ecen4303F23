magic
tech scmos
timestamp 1071163401
<< nwell >>
rect -8 68 184 105
<< ntransistor >>
rect 8 6 10 26
rect 14 6 16 26
rect 24 6 26 26
rect 30 6 32 26
rect 47 6 49 16
rect 55 6 57 16
rect 63 6 65 16
rect 79 6 81 16
rect 87 6 89 16
rect 103 6 105 16
rect 111 6 113 16
rect 128 6 130 26
rect 134 6 136 26
rect 144 6 146 26
rect 150 6 152 26
rect 167 6 169 16
<< ptransistor >>
rect 7 74 9 94
rect 15 74 17 94
rect 23 74 25 94
rect 31 74 33 94
rect 47 84 49 94
rect 55 84 57 94
rect 63 74 65 94
rect 79 74 81 94
rect 87 74 89 94
rect 103 84 105 94
rect 111 84 113 94
rect 127 74 129 94
rect 135 74 137 94
rect 143 74 145 94
rect 151 74 153 94
rect 167 74 169 94
<< ndiffusion >>
rect 6 6 8 26
rect 10 6 14 26
rect 16 6 18 26
rect 22 6 24 26
rect 26 6 30 26
rect 32 6 34 26
rect 46 6 47 16
rect 49 6 50 16
rect 54 6 55 16
rect 57 6 58 16
rect 62 6 63 16
rect 65 6 66 16
rect 78 6 79 16
rect 81 6 82 16
rect 86 6 87 16
rect 89 6 90 16
rect 102 6 103 16
rect 105 6 106 16
rect 110 6 111 16
rect 113 6 114 16
rect 126 6 128 26
rect 130 6 134 26
rect 136 6 138 26
rect 142 6 144 26
rect 146 6 150 26
rect 152 6 154 26
rect 166 6 167 16
rect 169 6 170 16
<< pdiffusion >>
rect 6 74 7 94
rect 9 74 10 94
rect 14 74 15 94
rect 17 74 18 94
rect 22 74 23 94
rect 25 74 26 94
rect 30 74 31 94
rect 33 74 34 94
rect 46 84 47 94
rect 49 84 50 94
rect 54 84 55 94
rect 57 84 58 94
rect 62 74 63 94
rect 65 74 66 94
rect 78 74 79 94
rect 81 74 82 94
rect 86 74 87 94
rect 89 74 90 94
rect 102 84 103 94
rect 105 84 106 94
rect 110 84 111 94
rect 113 84 114 94
rect 126 74 127 94
rect 129 74 130 94
rect 134 74 135 94
rect 137 74 138 94
rect 142 74 143 94
rect 145 74 146 94
rect 150 74 151 94
rect 153 74 154 94
rect 166 74 167 94
rect 169 74 170 94
<< ndcontact >>
rect 2 6 6 26
rect 18 6 22 26
rect 34 6 38 26
rect 42 6 46 16
rect 50 6 54 16
rect 58 6 62 16
rect 66 6 70 16
rect 74 6 78 16
rect 82 6 86 16
rect 90 6 94 16
rect 98 6 102 16
rect 106 6 110 16
rect 114 6 118 16
rect 122 6 126 26
rect 138 6 142 26
rect 154 6 158 26
rect 162 6 166 16
rect 170 6 174 16
<< pdcontact >>
rect 2 74 6 94
rect 10 74 14 94
rect 18 74 22 94
rect 26 74 30 94
rect 34 74 38 94
rect 42 84 46 94
rect 50 84 54 94
rect 58 74 62 94
rect 66 74 70 94
rect 74 74 78 94
rect 82 74 86 94
rect 90 74 94 94
rect 98 84 102 94
rect 106 84 110 94
rect 114 84 118 94
rect 122 74 126 94
rect 130 74 134 94
rect 138 74 142 94
rect 146 74 150 94
rect 154 74 158 94
rect 162 74 166 94
rect 170 74 174 94
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
rect 46 -2 50 2
rect 62 -2 66 2
rect 78 -2 82 2
rect 94 -2 98 2
rect 110 -2 114 2
rect 126 -2 130 2
rect 142 -2 146 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
rect 46 98 50 102
rect 62 98 66 102
rect 78 98 82 102
rect 94 98 98 102
rect 110 98 114 102
rect 126 98 130 102
rect 142 98 146 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 31 94 33 96
rect 47 94 49 96
rect 55 94 57 96
rect 63 94 65 96
rect 79 94 81 96
rect 87 94 89 96
rect 103 94 105 96
rect 111 94 113 96
rect 127 94 129 96
rect 135 94 137 96
rect 143 94 145 96
rect 151 94 153 96
rect 167 94 169 96
rect 7 73 9 74
rect 4 71 9 73
rect 4 48 6 71
rect 15 65 17 74
rect 14 61 17 65
rect 15 56 17 61
rect 23 64 25 74
rect 31 71 33 74
rect 47 73 49 84
rect 47 71 51 73
rect 31 69 35 71
rect 15 54 19 56
rect 4 44 9 48
rect 4 29 6 44
rect 17 33 19 54
rect 18 29 19 33
rect 23 29 25 60
rect 33 51 35 69
rect 31 49 35 51
rect 31 30 33 49
rect 49 42 51 71
rect 55 67 57 84
rect 103 83 105 84
rect 101 81 105 83
rect 63 73 65 74
rect 63 71 75 73
rect 55 63 65 67
rect 57 34 59 63
rect 73 59 75 71
rect 79 70 81 74
rect 87 73 89 74
rect 4 27 10 29
rect 8 26 10 27
rect 14 26 16 29
rect 23 27 26 29
rect 24 26 26 27
rect 30 28 33 30
rect 47 32 59 34
rect 63 57 75 59
rect 78 68 81 70
rect 84 71 89 73
rect 63 33 65 57
rect 78 42 80 68
rect 84 59 86 71
rect 101 67 103 81
rect 111 71 113 84
rect 94 63 103 67
rect 84 57 88 59
rect 30 26 32 28
rect 47 16 49 32
rect 63 29 66 33
rect 55 16 57 23
rect 63 16 65 29
rect 78 19 80 38
rect 86 27 88 57
rect 101 47 103 63
rect 100 45 103 47
rect 106 69 113 71
rect 96 31 97 35
rect 100 33 102 45
rect 106 41 110 69
rect 127 60 129 74
rect 135 73 137 74
rect 114 58 129 60
rect 133 71 137 73
rect 114 38 116 58
rect 133 54 135 71
rect 143 56 145 74
rect 129 52 135 54
rect 138 54 145 56
rect 151 54 153 74
rect 129 46 131 52
rect 126 42 131 46
rect 138 42 140 54
rect 114 36 120 38
rect 100 31 115 33
rect 95 27 97 31
rect 95 25 105 27
rect 78 17 81 19
rect 79 16 81 17
rect 87 16 89 23
rect 103 16 105 25
rect 113 19 115 31
rect 118 29 120 36
rect 129 34 131 42
rect 139 38 140 42
rect 138 34 140 38
rect 144 50 149 51
rect 144 49 153 50
rect 144 34 146 49
rect 167 42 169 74
rect 154 38 169 42
rect 129 32 135 34
rect 138 32 141 34
rect 144 32 152 34
rect 133 29 135 32
rect 139 29 141 32
rect 118 27 130 29
rect 133 27 136 29
rect 139 27 146 29
rect 128 26 130 27
rect 134 26 136 27
rect 144 26 146 27
rect 150 26 152 32
rect 111 17 115 19
rect 111 16 113 17
rect 167 16 169 38
rect 8 4 10 6
rect 14 4 16 6
rect 24 4 26 6
rect 30 4 32 6
rect 47 4 49 6
rect 55 4 57 6
rect 63 4 65 6
rect 79 4 81 6
rect 87 4 89 6
rect 103 4 105 6
rect 111 4 113 6
rect 128 4 130 6
rect 134 4 136 6
rect 144 4 146 6
rect 150 4 152 6
rect 167 4 169 6
<< polycontact >>
rect 10 61 14 65
rect 23 60 27 64
rect 9 44 13 48
rect 14 29 18 33
rect 35 51 39 55
rect 65 63 69 67
rect 49 38 53 42
rect 90 63 94 67
rect 78 38 82 42
rect 66 29 70 33
rect 55 23 59 27
rect 74 23 78 27
rect 92 31 96 35
rect 123 67 127 71
rect 106 37 110 41
rect 139 63 143 67
rect 122 42 126 46
rect 86 23 90 27
rect 105 23 109 27
rect 135 38 139 42
rect 149 50 153 54
rect 150 38 154 42
<< metal1 >>
rect -2 102 178 103
rect 2 98 14 102
rect 18 98 30 102
rect 34 98 46 102
rect 50 98 62 102
rect 66 98 78 102
rect 82 98 94 102
rect 98 98 110 102
rect 114 98 126 102
rect 130 98 142 102
rect 146 98 178 102
rect -2 97 178 98
rect 2 94 6 97
rect 18 94 22 97
rect 34 94 38 97
rect 66 94 70 97
rect 82 94 86 97
rect 122 94 126 97
rect 138 94 142 97
rect 154 94 158 97
rect 170 94 174 97
rect 9 74 10 77
rect 9 71 12 74
rect 26 71 30 74
rect 2 68 12 71
rect 2 40 6 68
rect 15 67 36 71
rect 90 67 94 70
rect 110 67 123 71
rect 130 67 134 74
rect 146 71 150 74
rect 146 68 159 71
rect 15 65 18 67
rect 14 61 18 65
rect 33 64 62 67
rect 27 61 30 64
rect 27 58 50 61
rect 59 60 62 64
rect 69 63 74 67
rect 130 63 139 67
rect 59 57 98 60
rect 156 60 159 68
rect 118 57 159 60
rect 18 54 22 57
rect 18 51 35 54
rect 39 51 149 54
rect 156 48 159 57
rect 162 55 166 74
rect 162 51 167 55
rect 13 46 126 48
rect 13 45 122 46
rect 34 43 38 45
rect 156 45 160 48
rect 2 36 42 40
rect 53 38 59 42
rect 82 38 90 42
rect 2 26 6 36
rect 18 29 29 33
rect 25 26 29 29
rect 55 27 59 38
rect 66 33 70 37
rect 78 31 92 34
rect 106 27 110 37
rect 139 38 150 42
rect 135 32 139 38
rect 157 35 160 45
rect 25 22 34 26
rect 59 23 74 26
rect 82 23 86 27
rect 109 23 110 27
rect 130 29 139 32
rect 154 32 160 35
rect 130 26 134 29
rect 154 26 158 32
rect 163 29 167 51
rect 126 22 134 26
rect 162 25 167 29
rect 162 16 166 25
rect 18 3 22 6
rect 66 3 70 6
rect 82 3 86 6
rect 138 3 142 6
rect 170 3 174 6
rect -2 2 178 3
rect 2 -2 14 2
rect 18 -2 30 2
rect 34 -2 46 2
rect 50 -2 62 2
rect 66 -2 78 2
rect 82 -2 94 2
rect 98 -2 110 2
rect 114 -2 126 2
rect 130 -2 142 2
rect 146 -2 178 2
rect -2 -3 178 -2
<< m2contact >>
rect 42 80 46 84
rect 50 80 54 84
rect 98 80 102 84
rect 106 80 110 84
rect 114 80 118 84
rect 58 70 62 74
rect 74 70 78 74
rect 90 70 94 74
rect 106 67 110 71
rect 50 57 54 61
rect 74 63 78 67
rect 98 57 102 61
rect 114 57 118 61
rect 42 36 46 40
rect 90 38 94 42
rect 74 30 78 34
rect 42 16 46 20
rect 50 16 54 20
rect 58 16 62 20
rect 74 16 78 20
rect 90 16 94 20
rect 98 16 102 20
rect 106 16 110 20
rect 114 16 118 20
<< metal2 >>
rect 42 40 46 80
rect 42 20 46 36
rect 50 61 54 80
rect 50 20 54 57
rect 58 20 62 70
rect 74 67 78 70
rect 74 34 78 63
rect 74 20 78 30
rect 90 42 94 70
rect 90 20 94 38
rect 98 61 102 80
rect 98 20 102 57
rect 106 71 110 80
rect 106 20 110 67
rect 114 61 118 80
rect 114 20 118 57
<< m1p >>
rect 162 63 166 67
rect 18 53 22 57
rect 34 43 38 47
rect 66 33 70 37
rect 82 23 86 27
<< labels >>
rlabel metal1 4 0 4 0 1 gnd
rlabel metal1 4 100 4 100 5 vdd
rlabel metal1 68 35 68 35 1 D
rlabel metal1 20 55 20 55 1 S
rlabel metal1 36 45 36 45 1 R
rlabel metal1 164 65 164 65 1 Q
rlabel metal1 84 25 84 25 1 CLK
<< end >>
